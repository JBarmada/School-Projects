module go_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [7:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin








		if(({row_reg, col_reg}>=14'b00000000000000) && ({row_reg, col_reg}<14'b00100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00100000000001) && ({row_reg, col_reg}<14'b00100000001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100000001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00100000001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00100000001100) && ({row_reg, col_reg}<14'b00100000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00100000010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00100000010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00100000010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00100000010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b00100000010100) && ({row_reg, col_reg}<14'b00100000010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b00100000010110) && ({row_reg, col_reg}<14'b00100000011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b00100000011000) && ({row_reg, col_reg}<14'b00100000011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00100000011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00100000011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100000011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00100000011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00100000011110) && ({row_reg, col_reg}<14'b00100001110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100001110000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00100001110001) && ({row_reg, col_reg}<14'b00100100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00100100001010) && ({row_reg, col_reg}<14'b00100100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100100001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00100100001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b00100100001111) && ({row_reg, col_reg}<14'b00100100010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b00100100010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b00100100010011) && ({row_reg, col_reg}<14'b00100100010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00100100010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b00100100010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b00100100010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b00100100011000) && ({row_reg, col_reg}<14'b00100100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00100100011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b00100100011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00100100011100) && ({row_reg, col_reg}<14'b00100100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100100011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00100100100000) && ({row_reg, col_reg}<14'b00100101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00100110000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00100110000001) && ({row_reg, col_reg}<14'b00100110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100110000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00100110000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00100110000101) && ({row_reg, col_reg}<14'b00100110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00100110000111)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b00100110001000) && ({row_reg, col_reg}<14'b00101000000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00101000000110) && ({row_reg, col_reg}<14'b00101000001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00101000001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00101000001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00101000001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b00101000001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101000010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00101000010001) && ({row_reg, col_reg}<14'b00101000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101000011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101000011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b00101000011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b00101000011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b00101000011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00101000011110) && ({row_reg, col_reg}<14'b00101001111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101001111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00101001111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00101001111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b00101001111101) && ({row_reg, col_reg}<14'b00101001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00101001111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b00101010000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00101010000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00101010000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101010000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101010000100) && ({row_reg, col_reg}<14'b00101010000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101010000111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00101010001000) && ({row_reg, col_reg}<14'b00101100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101100001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00101100001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b00101100001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b00101100001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b00101100001110) && ({row_reg, col_reg}<14'b00101100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101100010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00101100010011) && ({row_reg, col_reg}<14'b00101100010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00101100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00101100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00101100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101100011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00101100011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00101100011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00101100011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00101100011111) && ({row_reg, col_reg}<14'b00101101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101101111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00101101111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00101101111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b00101101111100) && ({row_reg, col_reg}<14'b00101101111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b00101101111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b00101110000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00101110000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b00101110000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00101110000100) && ({row_reg, col_reg}<14'b00101110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00101110000110)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b00101110000111) && ({row_reg, col_reg}<14'b00110000000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00110000000011) && ({row_reg, col_reg}<14'b00110000001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110000001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110000001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00110000001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00110000001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b00110000001100) && ({row_reg, col_reg}<14'b00110000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110000001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110000001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00110000010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b00110000010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b00110000010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b00110000010011) && ({row_reg, col_reg}<14'b00110000010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00110000010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b00110000010110) && ({row_reg, col_reg}<14'b00110000011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b00110000011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00110000011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b00110000011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110000011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00110000011100) && ({row_reg, col_reg}<14'b00110000011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00110000011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b00110000011111) && ({row_reg, col_reg}<14'b00110001110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110001110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00110001110011) && ({row_reg, col_reg}<14'b00110001111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110001111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00110001111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b00110001111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110001111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110001111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00110001111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00110001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110010000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00110010000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b00110010000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00110010000100)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=14'b00110010000101) && ({row_reg, col_reg}<14'b00110100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00110100000011) && ({row_reg, col_reg}<14'b00110100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110100001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00110100001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b00110100001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b00110100001011) && ({row_reg, col_reg}<14'b00110100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110100001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00110100001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b00110100001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b00110100010000) && ({row_reg, col_reg}<14'b00110100010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00110100010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110100010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110100010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b00110100010101) && ({row_reg, col_reg}<14'b00110100010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110100010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00110100011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00110100011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00110100011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b00110100011011) && ({row_reg, col_reg}<14'b00110100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00110100011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b00110100011110) && ({row_reg, col_reg}<14'b00110101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00110101110001) && ({row_reg, col_reg}<14'b00110101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00110101110011) && ({row_reg, col_reg}<14'b00110101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110101111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b00110101111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b00110101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b00110101111011) && ({row_reg, col_reg}<14'b00110101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110110000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00110110000011) && ({row_reg, col_reg}<14'b00110110000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b00110110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00110110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00110110000111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00110110001000) && ({row_reg, col_reg}<14'b00111000000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111000000011) && ({row_reg, col_reg}<14'b00111000000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111000000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111000000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111000001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b00111000001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00111000001010) && ({row_reg, col_reg}<14'b00111000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111000001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00111000001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00111000001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b00111000001111) && ({row_reg, col_reg}<14'b00111000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111000010001) && ({row_reg, col_reg}<14'b00111000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111000011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00111000011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00111000011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111000011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00111000011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111000011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111000011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111000100000) && ({row_reg, col_reg}<14'b00111001110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111001110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111001110011) && ({row_reg, col_reg}<14'b00111001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111001110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111001110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111001111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b00111001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b00111001111010) && ({row_reg, col_reg}<14'b00111001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00111001111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b00111001111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b00111001111110) && ({row_reg, col_reg}<14'b00111010000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b00111010000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b00111010000001) && ({row_reg, col_reg}<14'b00111010000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111010000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00111010000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b00111010000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b00111010000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b00111010000111) && ({row_reg, col_reg}<14'b00111100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111100000011) && ({row_reg, col_reg}<14'b00111100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111100000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b00111100000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00111100001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b00111100001001) && ({row_reg, col_reg}<14'b00111100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111100001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b00111100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00111100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b00111100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b00111100010000) && ({row_reg, col_reg}<14'b00111100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00111100010011) && ({row_reg, col_reg}<14'b00111100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111100010101) && ({row_reg, col_reg}<14'b00111100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00111100011000) && ({row_reg, col_reg}<14'b00111100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111100011010) && ({row_reg, col_reg}<14'b00111100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b00111100011100) && ({row_reg, col_reg}<14'b00111100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b00111100011110) && ({row_reg, col_reg}<14'b00111101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111101110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b00111101110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b00111101111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b00111101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00111101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111101111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b00111101111100) && ({row_reg, col_reg}<14'b00111101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b00111101111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b00111101111111) && ({row_reg, col_reg}<14'b00111110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00111110000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b00111110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b00111110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b00111110000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b00111110000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b00111110000110)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=14'b00111110000111) && ({row_reg, col_reg}<14'b01000000000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000000000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01000000000010) && ({row_reg, col_reg}<14'b01000000000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000000000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01000000000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01000000000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01000000001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000000001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000000001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01000000001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01000000001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01000000001101) && ({row_reg, col_reg}<14'b01000001110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000001110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01000001110010) && ({row_reg, col_reg}<14'b01000001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01000001110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01000001111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000001111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000001111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000001111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01000001111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01000001111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01000001111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000010000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000010000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01000010000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b01000010000011) && ({row_reg, col_reg}<14'b01000010000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000010000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01000010000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01000010000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000010001000) && ({row_reg, col_reg}<14'b01000010011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000010011001) && ({row_reg, col_reg}<14'b01000010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000010100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000010100011) && ({row_reg, col_reg}<14'b01000010100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000010100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000010101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01000010101001) && ({row_reg, col_reg}<14'b01000010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000010101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000010101101) && ({row_reg, col_reg}<14'b01000010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000010110001) && ({row_reg, col_reg}<14'b01000010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000011000011) && ({row_reg, col_reg}<14'b01000011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000011000101)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b01000011000110) && ({row_reg, col_reg}<14'b01000100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000100000010) && ({row_reg, col_reg}<14'b01000100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000100000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01000100000110) && ({row_reg, col_reg}<14'b01000100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01000100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000100001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01000100001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000100001101) && ({row_reg, col_reg}<14'b01000101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01000101011011) && ({row_reg, col_reg}<14'b01000101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000101011110) && ({row_reg, col_reg}<14'b01000101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000101110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01000101110010) && ({row_reg, col_reg}<14'b01000101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000101110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01000101110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01000101111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000101111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01000101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01000101111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01000101111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01000101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000101111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01000110000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01000110000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000110000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01000110000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01000110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01000110001000) && ({row_reg, col_reg}<14'b01000110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000110100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000110100010) && ({row_reg, col_reg}<14'b01000110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000110100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000110100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01000110101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01000110101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01000110101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01000110101100) && ({row_reg, col_reg}<14'b01000110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000110101110) && ({row_reg, col_reg}<14'b01000110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000110110100) && ({row_reg, col_reg}<14'b01000110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000110110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01000110110111) && ({row_reg, col_reg}<14'b01000110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01000110111011) && ({row_reg, col_reg}<14'b01000111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01000111000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}==14'b01000111000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01001000000000) && ({row_reg, col_reg}<14'b01001000000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001000000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001000000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001000000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01001000000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01001000001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001000001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01001000001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01001000001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01001000001100) && ({row_reg, col_reg}<14'b01001001011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001001011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001001011101) && ({row_reg, col_reg}<14'b01001001110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001001110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01001001110010) && ({row_reg, col_reg}<14'b01001001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001001110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001001110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01001001110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b01001001111000) && ({row_reg, col_reg}<14'b01001001111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01001001111010) && ({row_reg, col_reg}<14'b01001001111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01001001111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01001001111101) && ({row_reg, col_reg}<14'b01001001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001001111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001010000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001010000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01001010000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01001010000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001010000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001010000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01001010000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b01001010001000) && ({row_reg, col_reg}<14'b01001010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01001010100000) && ({row_reg, col_reg}<14'b01001010100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001010100010) && ({row_reg, col_reg}<14'b01001010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001010101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01001010110000) && ({row_reg, col_reg}<14'b01001010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01001010110010) && ({row_reg, col_reg}<14'b01001010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001010110100) && ({row_reg, col_reg}<14'b01001010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001010111101) && ({row_reg, col_reg}<14'b01001011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001011000001) && ({row_reg, col_reg}<14'b01001011000111)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==14'b01001011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01001100000000) && ({row_reg, col_reg}<14'b01001100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001100000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01001100000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01001100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001100001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001100001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01001100001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01001100001011) && ({row_reg, col_reg}<14'b01001101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001101110010) && ({row_reg, col_reg}<14'b01001101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001101110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001101110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01001101110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01001101111000) && ({row_reg, col_reg}<14'b01001101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001101111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01001101111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b01001101111100) && ({row_reg, col_reg}<14'b01001101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01001101111111) && ({row_reg, col_reg}<14'b01001110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001110000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01001110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01001110000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001110000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01001110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01001110001000) && ({row_reg, col_reg}<14'b01001110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001110010000) && ({row_reg, col_reg}<14'b01001110011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01001110011010) && ({row_reg, col_reg}<14'b01001110011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001110011100) && ({row_reg, col_reg}<14'b01001110011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001110100000) && ({row_reg, col_reg}<14'b01001110100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001110100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01001110100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01001110100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01001110101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01001110101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01001110101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01001110101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01001110101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01001110101101) && ({row_reg, col_reg}<14'b01001110110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001110110011) && ({row_reg, col_reg}<14'b01001110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001110110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01001110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001110111000) && ({row_reg, col_reg}<14'b01001111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01001111000001) && ({row_reg, col_reg}<14'b01001111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01001111000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01001111000100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01001111000101) && ({row_reg, col_reg}<14'b01010000000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010000000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01010000000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01010000000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010000001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01010000001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01010000001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010000001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010000001101) && ({row_reg, col_reg}<14'b01010000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010000001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010000010000) && ({row_reg, col_reg}<14'b01010001011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010001011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010001011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010001011010) && ({row_reg, col_reg}<14'b01010001011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010001011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010001100000) && ({row_reg, col_reg}<14'b01010001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010001110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010001110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01010001110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010001111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010001111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010001111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01010001111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01010001111100) && ({row_reg, col_reg}<14'b01010010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010010000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01010010000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010010000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01010010000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01010010000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01010010000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010010000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010010000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01010010001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010010001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010010001010) && ({row_reg, col_reg}<14'b01010010010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010010011000) && ({row_reg, col_reg}<14'b01010010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010010100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010010100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010010100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01010010100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01010010100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01010010101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01010010101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01010010101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01010010101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01010010101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01010010101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01010010101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01010010101111) && ({row_reg, col_reg}<14'b01010010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010010110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010010110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01010010110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b01010010111000) && ({row_reg, col_reg}<14'b01010010111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010010111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010010111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010010111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01010010111101) && ({row_reg, col_reg}<14'b01010010111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010010111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010011000000)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01010011000001) && ({row_reg, col_reg}<14'b01010100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010100000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01010100000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010100001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01010100001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01010100001010) && ({row_reg, col_reg}<14'b01010100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010100001101) && ({row_reg, col_reg}<14'b01010101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010101110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010101110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01010101110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010101111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010101111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01010101111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010101111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010101111110) && ({row_reg, col_reg}<14'b01010110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010110000001) && ({row_reg, col_reg}<14'b01010110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01010110000011) && ({row_reg, col_reg}<14'b01010110000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01010110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010110000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01010110001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01010110001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010110001010) && ({row_reg, col_reg}<14'b01010110001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01010110001101) && ({row_reg, col_reg}<14'b01010110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010110010001) && ({row_reg, col_reg}<14'b01010110011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010110011001) && ({row_reg, col_reg}<14'b01010110011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01010110011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01010110011100) && ({row_reg, col_reg}<14'b01010110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010110100001) && ({row_reg, col_reg}<14'b01010110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01010110100100) && ({row_reg, col_reg}<14'b01010110100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01010110100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01010110100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01010110101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01010110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010110101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01010110101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01010110101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01010110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01010110110001) && ({row_reg, col_reg}<14'b01010110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01010110110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01010110110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01010110110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01010110111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01010110111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01010110111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01010110111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01010110111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b01010110111101) && ({row_reg, col_reg}<14'b01010111000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01010111000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01010111000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01010111000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01010111000011) && ({row_reg, col_reg}<14'b01010111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01010111000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01010111000111) && ({row_reg, col_reg}<14'b01011000000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011000000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011000000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01011000000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011000001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01011000001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011000001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01011000001100) && ({row_reg, col_reg}<14'b01011001011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011001011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011001011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011001011101) && ({row_reg, col_reg}<14'b01011001011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01011001011111) && ({row_reg, col_reg}<14'b01011001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011001110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011001110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011001110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01011001110111) && ({row_reg, col_reg}<14'b01011001111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011001111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011001111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01011001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011001111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011001111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01011001111110) && ({row_reg, col_reg}<14'b01011010000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011010000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011010000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01011010000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011010000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011010000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01011010001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01011010001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011010001010) && ({row_reg, col_reg}<14'b01011010001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011010001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011010001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011010001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011010001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011010010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011010010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01011010010010) && ({row_reg, col_reg}<14'b01011010011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011010011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01011010011001) && ({row_reg, col_reg}<14'b01011010011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01011010011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011010011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011010011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01011010011111) && ({row_reg, col_reg}<14'b01011010100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011010100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011010100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01011010100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01011010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011010100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01011010100110) && ({row_reg, col_reg}<14'b01011010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011010101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01011010101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01011010101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01011010101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01011010101110) && ({row_reg, col_reg}<14'b01011010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01011010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011010110001) && ({row_reg, col_reg}<14'b01011010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011010110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011010110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01011010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011010111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01011010111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01011010111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011010111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011010111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011011000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01011011000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01011011000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01011011000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011011000100) && ({row_reg, col_reg}<14'b01011011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011011000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01011011000111) && ({row_reg, col_reg}<14'b01011100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01011100000010) && ({row_reg, col_reg}<14'b01011100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011100000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01011100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011100000111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011100001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01011100001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011100001100) && ({row_reg, col_reg}<14'b01011100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011100001111) && ({row_reg, col_reg}<14'b01011101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011101011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01011101011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011101011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011101011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011101011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011101011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01011101100000) && ({row_reg, col_reg}<14'b01011101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011101110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011101110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01011101110111) && ({row_reg, col_reg}<14'b01011101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011101111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01011101111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b01011101111011) && ({row_reg, col_reg}<14'b01011101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011101111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011101111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01011110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011110000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01011110000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01011110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01011110001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01011110001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011110001010) && ({row_reg, col_reg}<14'b01011110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01011110001101) && ({row_reg, col_reg}<14'b01011110010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01011110010000) && ({row_reg, col_reg}<14'b01011110010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011110010010) && ({row_reg, col_reg}<14'b01011110011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01011110011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01011110011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01011110011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011110011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01011110011101) && ({row_reg, col_reg}<14'b01011110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01011110100010) && ({row_reg, col_reg}<14'b01011110100100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01011110100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011110100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011110100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01011110101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01011110101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01011110101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01011110101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01011110101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01011110101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01011110101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01011110110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011110110001) && ({row_reg, col_reg}<14'b01011110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011110110101) && ({row_reg, col_reg}<14'b01011110110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01011110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01011110111010) && ({row_reg, col_reg}<14'b01011110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011110111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01011110111110) && ({row_reg, col_reg}<14'b01011111000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01011111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011111000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01011111000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01011111000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01011111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01011111000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01011111000110)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b01011111000111) && ({row_reg, col_reg}<14'b01100000000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100000000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100000000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100000000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100000000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100000001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100000001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100000001101) && ({row_reg, col_reg}<14'b01100000010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100000010010) && ({row_reg, col_reg}<14'b01100000010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100000010111) && ({row_reg, col_reg}<14'b01100000011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01100000011010) && ({row_reg, col_reg}<14'b01100000011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100000011100) && ({row_reg, col_reg}<14'b01100000100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100000100011) && ({row_reg, col_reg}<14'b01100000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100000100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01100000100111) && ({row_reg, col_reg}<14'b01100000110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01100000110100) && ({row_reg, col_reg}<14'b01100000110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100000110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100000111001) && ({row_reg, col_reg}<14'b01100000111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100000111100) && ({row_reg, col_reg}<14'b01100000111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100000111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100001000000) && ({row_reg, col_reg}<14'b01100001000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100001000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01100001000011) && ({row_reg, col_reg}<14'b01100001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100001001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100001001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100001001100) && ({row_reg, col_reg}<14'b01100001010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100001010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100001010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01100001010100) && ({row_reg, col_reg}<14'b01100001011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100001011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01100001011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01100001011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b01100001011011) && ({row_reg, col_reg}<14'b01100001011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100001011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b01100001011110) && ({row_reg, col_reg}<14'b01100001100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100001100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100001100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100001100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01100001100011) && ({row_reg, col_reg}<14'b01100001100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100001100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100001100110) && ({row_reg, col_reg}<14'b01100001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100001110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100001110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01100001110111) && ({row_reg, col_reg}<14'b01100001111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100001111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100001111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100001111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100001111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100001111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100010000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100010000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100010000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100010000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100010000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100010001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100010001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01100010001010) && ({row_reg, col_reg}<14'b01100010001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100010001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100010001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100010001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100010010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100010010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100010010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01100010010011) && ({row_reg, col_reg}<14'b01100010010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100010010101) && ({row_reg, col_reg}<14'b01100010010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100010011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100010011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100010011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100010011110) && ({row_reg, col_reg}<14'b01100010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100010100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b01100010100011) && ({row_reg, col_reg}<14'b01100010100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100010100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100010100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100010101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100010101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01100010101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100010101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100010101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01100010110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01100010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100010110010) && ({row_reg, col_reg}<14'b01100010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100010110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100010110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b01100010110111) && ({row_reg, col_reg}<14'b01100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100010111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100010111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100010111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01100010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100010111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100010111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100011000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100011000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01100011000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b01100011000100) && ({row_reg, col_reg}<14'b01100011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100011000110)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b01100011000111) && ({row_reg, col_reg}<14'b01100100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100100000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100100001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100100001100) && ({row_reg, col_reg}<14'b01100100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01100100010101) && ({row_reg, col_reg}<14'b01100100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100100010111) && ({row_reg, col_reg}<14'b01100100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100100100000) && ({row_reg, col_reg}<14'b01100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100100100110) && ({row_reg, col_reg}<14'b01100100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01100100101100) && ({row_reg, col_reg}<14'b01100100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100100101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100100110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100100110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100100110011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b01100100110100) && ({row_reg, col_reg}<14'b01100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100100111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100100111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01100100111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100101000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100101000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100101000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100101001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100101001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01100101001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100101001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01100101001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01100101001110) && ({row_reg, col_reg}<14'b01100101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100101010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100101010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01100101011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100101011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100101011011) && ({row_reg, col_reg}<14'b01100101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100101011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100101011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100101100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100101100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100101100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100101100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b01100101100100) && ({row_reg, col_reg}<14'b01100101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01100101101000) && ({row_reg, col_reg}<14'b01100101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100101110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100101110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01100101110111) && ({row_reg, col_reg}<14'b01100101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100101111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01100101111110) && ({row_reg, col_reg}<14'b01100110000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100110000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100110000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100110000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100110000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100110001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100110001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100110001010) && ({row_reg, col_reg}<14'b01100110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01100110001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100110001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100110001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100110010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100110010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01100110010010) && ({row_reg, col_reg}<14'b01100110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100110010101) && ({row_reg, col_reg}<14'b01100110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100110011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100110011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100110011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01100110011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100110011110) && ({row_reg, col_reg}<14'b01100110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100110100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100110100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100110100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100110100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100110100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100110101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100110101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100110101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01100110101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100110101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100110101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100110101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01100110110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01100110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01100110110010) && ({row_reg, col_reg}<14'b01100110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01100110110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100110110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01100110111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01100110111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01100110111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01100110111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01100110111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100110111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01100111000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01100111000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01100111000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01100111000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b01100111000100) && ({row_reg, col_reg}<14'b01100111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100111000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01100111000111) && ({row_reg, col_reg}<14'b01101000000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101000000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101000000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101000000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01101000000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101000000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101000001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101000001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101000001100) && ({row_reg, col_reg}<14'b01101000010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101000010001) && ({row_reg, col_reg}<14'b01101000010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101000010101) && ({row_reg, col_reg}<14'b01101000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101000100101) && ({row_reg, col_reg}<14'b01101000101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101000101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101000101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01101000101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101000101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101000101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101000101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01101000110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01101000110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101000110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101000110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101000110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101000110101) && ({row_reg, col_reg}<14'b01101000110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101000111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101000111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101000111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101000111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101000111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101000111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101000111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01101001000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101001000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101001000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101001000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101001000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101001000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001000111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101001001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101001001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101001001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101001001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101001001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101001001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101001001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01101001001111) && ({row_reg, col_reg}<14'b01101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101001010010) && ({row_reg, col_reg}<14'b01101001010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101001010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101001010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01101001011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101001011001) && ({row_reg, col_reg}<14'b01101001011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101001011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101001011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101001011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101001011111) && ({row_reg, col_reg}<14'b01101001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101001100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101001100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01101001100100) && ({row_reg, col_reg}<14'b01101001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101001101000) && ({row_reg, col_reg}<14'b01101001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01101001110111) && ({row_reg, col_reg}<14'b01101001111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101001111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101001111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101001111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101001111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01101001111110) && ({row_reg, col_reg}<14'b01101010000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101010000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101010000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101010000010) && ({row_reg, col_reg}<14'b01101010000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01101010000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101010000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101010001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01101010001001) && ({row_reg, col_reg}<14'b01101010001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101010001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101010001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101010001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101010010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101010010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101010010101) && ({row_reg, col_reg}<14'b01101010010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101010011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101010011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101010011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01101010011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01101010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101010011110) && ({row_reg, col_reg}<14'b01101010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101010100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b01101010100010) && ({row_reg, col_reg}<14'b01101010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101010101001) && ({row_reg, col_reg}<14'b01101010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101010101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101010110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01101010110001) && ({row_reg, col_reg}<14'b01101010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101010110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101010110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01101010111000) && ({row_reg, col_reg}<14'b01101010111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101010111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101010111101) && ({row_reg, col_reg}<14'b01101011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101011000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01101011000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101011000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101011000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01101011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101011000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01101011000111) && ({row_reg, col_reg}<14'b01101100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101100000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101100000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01101100000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101100000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101100001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101100001010) && ({row_reg, col_reg}<14'b01101100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101100010001) && ({row_reg, col_reg}<14'b01101100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101100011010) && ({row_reg, col_reg}<14'b01101100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01101100011100) && ({row_reg, col_reg}<14'b01101100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101100011110) && ({row_reg, col_reg}<14'b01101100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101100100010) && ({row_reg, col_reg}<14'b01101100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101100100101) && ({row_reg, col_reg}<14'b01101100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101100101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101100101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01101100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01101100101111) && ({row_reg, col_reg}<14'b01101100110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101100110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101100110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101100110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101100110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01101100110111) && ({row_reg, col_reg}<14'b01101100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101100111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101100111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101100111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101100111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01101100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101101000010) && ({row_reg, col_reg}<14'b01101101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101101000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101101000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101101001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b01101101001001) && ({row_reg, col_reg}<14'b01101101001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101101001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01101101001111) && ({row_reg, col_reg}<14'b01101101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101101010010) && ({row_reg, col_reg}<14'b01101101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01101101010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101101010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01101101010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01101101011000) && ({row_reg, col_reg}<14'b01101101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01101101011011) && ({row_reg, col_reg}<14'b01101101011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101101011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01101101011111) && ({row_reg, col_reg}<14'b01101101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101101100110) && ({row_reg, col_reg}<14'b01101101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101101110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01101101110111) && ({row_reg, col_reg}<14'b01101101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101101111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101110000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101110000010) && ({row_reg, col_reg}<14'b01101110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01101110000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101110001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01101110001001) && ({row_reg, col_reg}<14'b01101110001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101110001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01101110010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01101110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01101110010011) && ({row_reg, col_reg}<14'b01101110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101110011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101110011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01101110011010) && ({row_reg, col_reg}<14'b01101110011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b01101110011100) && ({row_reg, col_reg}<14'b01101110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01101110100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101110100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01101110100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01101110100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101110100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b01101110101000) && ({row_reg, col_reg}<14'b01101110110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01101110110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01101110110001) && ({row_reg, col_reg}<14'b01101110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101110110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101110110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101110111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01101110111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01101110111010) && ({row_reg, col_reg}<14'b01101110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01101110111101) && ({row_reg, col_reg}<14'b01101110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01101110111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01101111000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01101111000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01101111000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01101111000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01101111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01101111000101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b01101111000110) && ({row_reg, col_reg}<14'b01110000000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110000000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01110000000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110000000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110000001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01110000001010) && ({row_reg, col_reg}<14'b01110000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110000001111) && ({row_reg, col_reg}<14'b01110000010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110000010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01110000011000) && ({row_reg, col_reg}<14'b01110000100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110000100100) && ({row_reg, col_reg}<14'b01110000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110000100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110000101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01110000101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01110000101010) && ({row_reg, col_reg}<14'b01110000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01110000101110) && ({row_reg, col_reg}<14'b01110000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110000110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110000110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110000110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01110000110110) && ({row_reg, col_reg}<14'b01110000111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110000111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110000111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110000111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110000111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110000111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110000111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110001000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110001000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110001000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110001000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110001000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110001000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110001000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110001001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110001001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110001001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110001001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01110001001100) && ({row_reg, col_reg}<14'b01110001001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110001001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110001010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110001010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110001010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110001010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01110001010111) && ({row_reg, col_reg}<14'b01110001011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110001011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01110001011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110001011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110001011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110001011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01110001011111) && ({row_reg, col_reg}<14'b01110001100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110001100001) && ({row_reg, col_reg}<14'b01110001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110001100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01110001100110) && ({row_reg, col_reg}<14'b01110001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01110001110111) && ({row_reg, col_reg}<14'b01110001111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01110001111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110001111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01110001111101) && ({row_reg, col_reg}<14'b01110010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01110010000001) && ({row_reg, col_reg}<14'b01110010000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110010000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110010000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110010000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110010001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110010001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110010001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110010001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110010001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01110010001111) && ({row_reg, col_reg}<14'b01110010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01110010010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01110010010011) && ({row_reg, col_reg}<14'b01110010010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110010010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110010011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110010011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110010011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110010011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01110010011100) && ({row_reg, col_reg}<14'b01110010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110010100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110010100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110010100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110010100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110010100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110010101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01110010101001) && ({row_reg, col_reg}<14'b01110010101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01110010101011) && ({row_reg, col_reg}<14'b01110010101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110010101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110010110001) && ({row_reg, col_reg}<14'b01110010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110010110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110010111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01110010111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01110010111010) && ({row_reg, col_reg}<14'b01110011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110011000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110011000010)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b01110011000011) && ({row_reg, col_reg}<14'b01110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110100000001) && ({row_reg, col_reg}<14'b01110100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01110100000011) && ({row_reg, col_reg}<14'b01110100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110100000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01110100000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110100001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01110100001010) && ({row_reg, col_reg}<14'b01110100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110100001111) && ({row_reg, col_reg}<14'b01110100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110100010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110100010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110100011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110100011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b01110100011010) && ({row_reg, col_reg}<14'b01110100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110100011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01110100011101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110100011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110100100001) && ({row_reg, col_reg}<14'b01110100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110100100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110100100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b01110100101000) && ({row_reg, col_reg}<14'b01110100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110100101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110100101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110100101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01110100110000) && ({row_reg, col_reg}<14'b01110100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110100110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01110100110101) && ({row_reg, col_reg}<14'b01110100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01110100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01110100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110100111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110101000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110101000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110101000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110101000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110101000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01110101000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110101000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110101001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01110101001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110101001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110101001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110101010010) && ({row_reg, col_reg}<14'b01110101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110101010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b01110101010110) && ({row_reg, col_reg}<14'b01110101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01110101011010) && ({row_reg, col_reg}<14'b01110101011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110101100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110101100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01110101100100) && ({row_reg, col_reg}<14'b01110101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110101100110) && ({row_reg, col_reg}<14'b01110101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110101110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01110101110111) && ({row_reg, col_reg}<14'b01110101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01110101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110101111101) && ({row_reg, col_reg}<14'b01110101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110110000000) && ({row_reg, col_reg}<14'b01110110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110110000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01110110000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110110001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01110110001001) && ({row_reg, col_reg}<14'b01110110001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01110110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110110001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110110001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01110110010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110110010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110110010100) && ({row_reg, col_reg}<14'b01110110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110110010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110110011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110110011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01110110011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01110110011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b01110110011100) && ({row_reg, col_reg}<14'b01110110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110110011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110110100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01110110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01110110100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01110110100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110110100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01110110101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01110110101010) && ({row_reg, col_reg}<14'b01110110110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01110110110011) && ({row_reg, col_reg}<14'b01110110110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110110110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01110110110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01110110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01110110111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01110110111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01110110111010) && ({row_reg, col_reg}<14'b01110111000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110111000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01110111000010) && ({row_reg, col_reg}<14'b01110111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01110111000110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}==14'b01110111000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111000000001) && ({row_reg, col_reg}<14'b01111000000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111000000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111000000110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111000000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111000001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111000001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01111000001010) && ({row_reg, col_reg}<14'b01111000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111000001100) && ({row_reg, col_reg}<14'b01111000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111000001111) && ({row_reg, col_reg}<14'b01111000010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111000010010) && ({row_reg, col_reg}<14'b01111000010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111000010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111000010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111000010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111000011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111000011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111000011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111000011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01111000011100) && ({row_reg, col_reg}<14'b01111000011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111000011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111000011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01111000100001) && ({row_reg, col_reg}<14'b01111000100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111000100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111000100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111000101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111000101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111000101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111000101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01111000101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111000101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111000110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111000110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111000110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01111000110101) && ({row_reg, col_reg}<14'b01111000110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111000111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111000111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01111000111011) && ({row_reg, col_reg}<14'b01111000111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111000111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111000111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111000111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01111001000000) && ({row_reg, col_reg}<14'b01111001000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111001000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111001000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111001000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111001000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111001001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111001001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111001001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111001001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01111001001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111001010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111001010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111001010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111001011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111001011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01111001011010) && ({row_reg, col_reg}<14'b01111001011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111001011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111001100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111001100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b01111001100010) && ({row_reg, col_reg}<14'b01111001100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111001100101) && ({row_reg, col_reg}<14'b01111001110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01111001110111) && ({row_reg, col_reg}<14'b01111001111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111001111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111001111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111001111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111010000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111010000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111010000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111010000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111010000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01111010000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111010001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111010001001) && ({row_reg, col_reg}<14'b01111010001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111010001100) && ({row_reg, col_reg}<14'b01111010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111010001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01111010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111010010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111010010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b01111010010100) && ({row_reg, col_reg}<14'b01111010010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111010010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111010011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111010011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111010011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111010011100) && ({row_reg, col_reg}<14'b01111010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111010011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111010100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111010100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111010100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111010100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111010100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111010101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111010101001) && ({row_reg, col_reg}<14'b01111010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111010110000) && ({row_reg, col_reg}<14'b01111010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111010110011) && ({row_reg, col_reg}<14'b01111010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01111010110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111010111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111010111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01111010111111) && ({row_reg, col_reg}<14'b01111011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111011000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111011000110)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=14'b01111011000111) && ({row_reg, col_reg}<14'b01111100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111100000001) && ({row_reg, col_reg}<14'b01111100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111100000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111100000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111100001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111100001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111100001100) && ({row_reg, col_reg}<14'b01111100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111100001111) && ({row_reg, col_reg}<14'b01111100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111100010010) && ({row_reg, col_reg}<14'b01111100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111100010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111100010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111100010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111100011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111100011010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111100011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111100011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111100100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b01111100100001) && ({row_reg, col_reg}<14'b01111100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111100101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111100101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111100101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111100110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111100110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111100110110) && ({row_reg, col_reg}<14'b01111100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111100111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01111100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111100111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111100111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111101000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01111101000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01111101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111101000110) && ({row_reg, col_reg}<14'b01111101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111101001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111101001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01111101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01111101001011) && ({row_reg, col_reg}<14'b01111101001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b01111101001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111101001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111101001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111101010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111101010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111101010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111101010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111101010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b01111101011000) && ({row_reg, col_reg}<14'b01111101100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111101100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111101100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111101100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01111101100011) && ({row_reg, col_reg}<14'b01111101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111101110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111101110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b01111101110111) && ({row_reg, col_reg}<14'b01111101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01111101111100) && ({row_reg, col_reg}<14'b01111101111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111101111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b01111110000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111110000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b01111110000010) && ({row_reg, col_reg}<14'b01111110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111110000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b01111110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111110000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b01111110001000) && ({row_reg, col_reg}<14'b01111110001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111110001100) && ({row_reg, col_reg}<14'b01111110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b01111110001110) && ({row_reg, col_reg}<14'b01111110010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b01111110010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b01111110010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01111110010100) && ({row_reg, col_reg}<14'b01111110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01111110010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111110011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b01111110011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b01111110011011) && ({row_reg, col_reg}<14'b01111110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111110011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b01111110100001) && ({row_reg, col_reg}<14'b01111110100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b01111110100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b01111110100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b01111110100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111110100111) && ({row_reg, col_reg}<14'b01111110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111110101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111110101101) && ({row_reg, col_reg}<14'b01111110110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111110110011) && ({row_reg, col_reg}<14'b01111110110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b01111110110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b01111110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111110111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b01111110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b01111110111100) && ({row_reg, col_reg}<14'b01111110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b01111110111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b01111111000001) && ({row_reg, col_reg}<14'b01111111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111111000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b01111111000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01111111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01111111000110)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b01111111000111) && ({row_reg, col_reg}<14'b10000000000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000000000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10000000000111) && ({row_reg, col_reg}<14'b10000000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000000001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000000001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000000001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000000001101) && ({row_reg, col_reg}<14'b10000000010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000000010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10000000010111) && ({row_reg, col_reg}<14'b10000000011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b10000000011001) && ({row_reg, col_reg}<14'b10000000011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000000011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000000011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b10000000011101) && ({row_reg, col_reg}<14'b10000000011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10000000011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b10000000100000) && ({row_reg, col_reg}<14'b10000000100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000000100010) && ({row_reg, col_reg}<14'b10000000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10000000100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000000100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000000101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000000101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000000101101) && ({row_reg, col_reg}<14'b10000000101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000000110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000000110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000000110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10000000110101) && ({row_reg, col_reg}<14'b10000000111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000000111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10000000111011) && ({row_reg, col_reg}<14'b10000000111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000000111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000000111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000000111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000001000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000001000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000001000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000001000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000001000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000001001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b10000001001001) && ({row_reg, col_reg}<14'b10000001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000001001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000001001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000001001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000001001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000001010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000001010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10000001010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000001010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000001010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000001011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000001011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10000001011010) && ({row_reg, col_reg}<14'b10000001011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000001100000) && ({row_reg, col_reg}<14'b10000001100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10000001100010) && ({row_reg, col_reg}<14'b10000001100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000001100100) && ({row_reg, col_reg}<14'b10000001110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000001110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000001110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000001110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b10000001110111) && ({row_reg, col_reg}<14'b10000001111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10000001111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10000001111011) && ({row_reg, col_reg}<14'b10000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000001111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000001111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10000001111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000010000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000010000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10000010000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000010000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000010000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000010000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000010001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10000010001001) && ({row_reg, col_reg}<14'b10000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000010001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10000010010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000010010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b10000010010100) && ({row_reg, col_reg}<14'b10000010010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000010010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000010011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000010011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10000010011011) && ({row_reg, col_reg}<14'b10000010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000010100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000010100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000010100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b10000010100100) && ({row_reg, col_reg}<14'b10000010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10000010101010) && ({row_reg, col_reg}<14'b10000010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000010101101) && ({row_reg, col_reg}<14'b10000010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10000010110011) && ({row_reg, col_reg}<14'b10000010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010110101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10000010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000010111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10000010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000010111011)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=14'b10000010111100) && ({row_reg, col_reg}<14'b10000100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000100000011) && ({row_reg, col_reg}<14'b10000100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000100000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000100000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000100001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000100001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000100001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000100001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000100001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10000100010000) && ({row_reg, col_reg}<14'b10000100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000100010011) && ({row_reg, col_reg}<14'b10000100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000100010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10000100011000) && ({row_reg, col_reg}<14'b10000100011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000100011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000100011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000100011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000100011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10000100011110) && ({row_reg, col_reg}<14'b10000100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000100100001) && ({row_reg, col_reg}<14'b10000100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000100100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10000100100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000100101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10000100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10000100101011) && ({row_reg, col_reg}<14'b10000100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10000100101110) && ({row_reg, col_reg}<14'b10000100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000100110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000100110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000100110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10000100110101) && ({row_reg, col_reg}<14'b10000100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000100111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10000100111011) && ({row_reg, col_reg}<14'b10000100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000100111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000101000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000101001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b10000101001001) && ({row_reg, col_reg}<14'b10000101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000101001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000101001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000101010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000101010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10000101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000101010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10000101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000101011001) && ({row_reg, col_reg}<14'b10000101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000101011101) && ({row_reg, col_reg}<14'b10000101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10000101110010) && ({row_reg, col_reg}<14'b10000101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000101110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10000101111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000101111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000110000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10000110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000110000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10000110000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10000110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000110001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10000110001001) && ({row_reg, col_reg}<14'b10000110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000110001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000110010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000110010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000110010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000110010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000110010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000110010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10000110011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10000110011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000110011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10000110011011) && ({row_reg, col_reg}<14'b10000110011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000110100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10000110100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000110100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000110100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000110100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000110100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10000110100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10000110100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000110101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10000110101010) && ({row_reg, col_reg}<14'b10000110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10000110110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10000110110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10000110110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10000110111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10000110111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10000110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10000110111100) && ({row_reg, col_reg}<14'b10000110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10000110111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10000110111111) && ({row_reg, col_reg}<14'b10001000000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001000000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001000000011) && ({row_reg, col_reg}<14'b10001000000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001000000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10001000000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10001000001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001000001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10001000001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b10001000001100) && ({row_reg, col_reg}<14'b10001000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001000001111) && ({row_reg, col_reg}<14'b10001000011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10001000011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001000011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001000011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10001000011110) && ({row_reg, col_reg}<14'b10001000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001000100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10001000100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001000100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001000101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10001000101010) && ({row_reg, col_reg}<14'b10001000101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001000101101) && ({row_reg, col_reg}<14'b10001000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10001000110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001000110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001000110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10001000110110) && ({row_reg, col_reg}<14'b10001000111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001000111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10001000111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10001000111011) && ({row_reg, col_reg}<14'b10001000111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001000111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10001000111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001001000000) && ({row_reg, col_reg}<14'b10001001000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001001000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001001000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001001000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001001000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001001000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10001001001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10001001001001) && ({row_reg, col_reg}<14'b10001001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001001001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001001001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001001001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001001001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10001001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10001001010000) && ({row_reg, col_reg}<14'b10001001010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001001010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001001010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10001001010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001001010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001001010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10001001010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10001001011000) && ({row_reg, col_reg}<14'b10001001011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10001001011011) && ({row_reg, col_reg}<14'b10001001011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001001011101) && ({row_reg, col_reg}<14'b10001001110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001001110001) && ({row_reg, col_reg}<14'b10001001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001001110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10001001110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001001110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001001111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001001111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001001111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10001001111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001001111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10001001111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001010000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001010000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001010000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001010000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001010000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001010000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10001010001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001010001001) && ({row_reg, col_reg}<14'b10001010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001010001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001010010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b10001010010001) && ({row_reg, col_reg}<14'b10001010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001010010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001010010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10001010010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001010010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10001010011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001010011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10001010011011) && ({row_reg, col_reg}<14'b10001010011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001010100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001010100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10001010100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b10001010100101) && ({row_reg, col_reg}<14'b10001010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10001010101000) && ({row_reg, col_reg}<14'b10001010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001010110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10001010110010) && ({row_reg, col_reg}<14'b10001010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001010110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001010110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10001010110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001010111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001010111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10001010111010) && ({row_reg, col_reg}<14'b10001010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001010111110)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10001010111111) && ({row_reg, col_reg}<14'b10001100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001100000010) && ({row_reg, col_reg}<14'b10001100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001100000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10001100001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001100001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001100001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10001100001101) && ({row_reg, col_reg}<14'b10001100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001100010001) && ({row_reg, col_reg}<14'b10001100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001100010100) && ({row_reg, col_reg}<14'b10001100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001100010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001100011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001100011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10001100011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10001100100000) && ({row_reg, col_reg}<14'b10001100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001100100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001100100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10001100101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001100101100) && ({row_reg, col_reg}<14'b10001100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10001100110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001100110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10001100110110) && ({row_reg, col_reg}<14'b10001100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10001100111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10001100111111) && ({row_reg, col_reg}<14'b10001101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001101000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10001101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001101000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10001101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10001101001001) && ({row_reg, col_reg}<14'b10001101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001101001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001101001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10001101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10001101010001) && ({row_reg, col_reg}<14'b10001101010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001101010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10001101010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001101010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001101011001) && ({row_reg, col_reg}<14'b10001101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10001101011111) && ({row_reg, col_reg}<14'b10001101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001101100010) && ({row_reg, col_reg}<14'b10001101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001101110001) && ({row_reg, col_reg}<14'b10001101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001101110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001101110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001101110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10001101111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10001101111100) && ({row_reg, col_reg}<14'b10001101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001101111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001110000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10001110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10001110000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b10001110001000) && ({row_reg, col_reg}<14'b10001110001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10001110001100) && ({row_reg, col_reg}<14'b10001110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001110010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001110010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10001110010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001110010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10001110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10001110010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001110011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001110011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10001110011010) && ({row_reg, col_reg}<14'b10001110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001110100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10001110100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001110100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10001110101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10001110101100) && ({row_reg, col_reg}<14'b10001110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10001110101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10001110110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10001110110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10001110110010) && ({row_reg, col_reg}<14'b10001110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10001110110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10001110110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10001110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10001110111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b10001110111010) && ({row_reg, col_reg}<14'b10001110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10001110111100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10001110111101) && ({row_reg, col_reg}<14'b10010000000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010000000010) && ({row_reg, col_reg}<14'b10010000000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10010000000101) && ({row_reg, col_reg}<14'b10010000000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010000001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010000001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010000001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010000001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10010000001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010000001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10010000001111) && ({row_reg, col_reg}<14'b10010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010000011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010000011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010000011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010000011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10010000011110) && ({row_reg, col_reg}<14'b10010000100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010000100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010000100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010000100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010000100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10010000101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10010000101010) && ({row_reg, col_reg}<14'b10010000101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010000101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10010000110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010000110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010000110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010000110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010000110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10010000110101) && ({row_reg, col_reg}<14'b10010000111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010000111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010000111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010000111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010000111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10010000111111) && ({row_reg, col_reg}<14'b10010001000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010001000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010001000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10010001001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10010001001001) && ({row_reg, col_reg}<14'b10010001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010001001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010001001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010001001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010001001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010001010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010001010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010001010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010001010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010001010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010001011001) && ({row_reg, col_reg}<14'b10010001011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010001100000) && ({row_reg, col_reg}<14'b10010001110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010001110001) && ({row_reg, col_reg}<14'b10010001110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010001110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010001110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010001111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010001111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010001111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010001111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010001111101) && ({row_reg, col_reg}<14'b10010001111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010001111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010010000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010010000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010010000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10010010000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10010010000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b10010010001000) && ({row_reg, col_reg}<14'b10010010001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010010010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10010010010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010010010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010010010011) && ({row_reg, col_reg}<14'b10010010010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010010010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010010011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010010011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010010011010) && ({row_reg, col_reg}<14'b10010010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010010011101) && ({row_reg, col_reg}<14'b10010010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010010100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010010100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010010100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010010100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10010010100111) && ({row_reg, col_reg}<14'b10010010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010010101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010010101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010010110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010010110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b10010010110010) && ({row_reg, col_reg}<14'b10010010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010010110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010010111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010010111100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10010010111101) && ({row_reg, col_reg}<14'b10010100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010100000101) && ({row_reg, col_reg}<14'b10010100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010100001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010100001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010100001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010100001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010100001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010100001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010100010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010100010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010100010011) && ({row_reg, col_reg}<14'b10010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010100011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010100011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010100011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010100011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010100011111) && ({row_reg, col_reg}<14'b10010100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010100100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010100100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010100101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10010100101010) && ({row_reg, col_reg}<14'b10010100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010100101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010100101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010100110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010100110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010100110111) && ({row_reg, col_reg}<14'b10010100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10010100111011) && ({row_reg, col_reg}<14'b10010100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10010100111111) && ({row_reg, col_reg}<14'b10010101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010101000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010101000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10010101001001) && ({row_reg, col_reg}<14'b10010101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010101001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10010101001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10010101001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010101001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010101001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010101010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010101010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010101010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010101010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10010101010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010101010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10010101011000) && ({row_reg, col_reg}<14'b10010101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10010101011011) && ({row_reg, col_reg}<14'b10010101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010101011101) && ({row_reg, col_reg}<14'b10010101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010101100100) && ({row_reg, col_reg}<14'b10010101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010101101000) && ({row_reg, col_reg}<14'b10010101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010101110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10010101110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010101110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010101111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10010101111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010101111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10010101111101) && ({row_reg, col_reg}<14'b10010110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010110000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010110000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010110000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10010110000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010110000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10010110001000) && ({row_reg, col_reg}<14'b10010110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010110010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010110010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10010110010011) && ({row_reg, col_reg}<14'b10010110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010110010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10010110011001) && ({row_reg, col_reg}<14'b10010110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010110011100) && ({row_reg, col_reg}<14'b10010110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010110011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010110100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10010110100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010110100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10010110100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10010110101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10010110101001) && ({row_reg, col_reg}<14'b10010110101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10010110101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010110101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10010110101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010110101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10010110110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10010110110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010110110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10010110110011) && ({row_reg, col_reg}<14'b10010110110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010110110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10010110110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10010110111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010110111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10010110111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10010110111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10010110111100)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b10010110111101) && ({row_reg, col_reg}<14'b10011000000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011000000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011000000100) && ({row_reg, col_reg}<14'b10011000001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011000001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011000001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011000001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011000001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011000001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011000010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b10011000010001) && ({row_reg, col_reg}<14'b10011000010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011000010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011000010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011000010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011000010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10011000011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10011000011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10011000011010) && ({row_reg, col_reg}<14'b10011000011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011000011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011000011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10011000011110) && ({row_reg, col_reg}<14'b10011000100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10011000100000) && ({row_reg, col_reg}<14'b10011000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011000100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011000100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011000100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011000100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011000101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011000101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011000101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011000101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011000101100) && ({row_reg, col_reg}<14'b10011000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10011000101110) && ({row_reg, col_reg}<14'b10011000110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011000110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10011000110001) && ({row_reg, col_reg}<14'b10011000110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011000110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011000110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011000110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10011000110110) && ({row_reg, col_reg}<14'b10011000111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011000111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011000111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10011000111011) && ({row_reg, col_reg}<14'b10011000111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011000111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10011000111111) && ({row_reg, col_reg}<14'b10011001000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011001000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011001000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011001001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011001001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011001001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011001001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011001001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011001010010) && ({row_reg, col_reg}<14'b10011001010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b10011001010101) && ({row_reg, col_reg}<14'b10011001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011001010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10011001011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011001011001) && ({row_reg, col_reg}<14'b10011001011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011001011101) && ({row_reg, col_reg}<14'b10011001100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011001100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011001100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011001100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011001100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011001100101) && ({row_reg, col_reg}<14'b10011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011001101000) && ({row_reg, col_reg}<14'b10011001110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011001110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011001111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011001111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011001111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011001111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011001111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10011001111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011001111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011001111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011010000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011010000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011010000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011010000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011010000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011010000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011010000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b10011010000111) && ({row_reg, col_reg}<14'b10011010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011010010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011010010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011010010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011010010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011010010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011010010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011010010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011010010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011010011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011010011001) && ({row_reg, col_reg}<14'b10011010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011010011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011010011100) && ({row_reg, col_reg}<14'b10011010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011010011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011010011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011010100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011010100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10011010100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011010100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011010100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011010100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10011010100111) && ({row_reg, col_reg}<14'b10011010101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b10011010101001) && ({row_reg, col_reg}<14'b10011010101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b10011010101011) && ({row_reg, col_reg}<14'b10011010101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011010101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011010101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011010110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011010110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011010110011) && ({row_reg, col_reg}<14'b10011010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011010110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10011010111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011010111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011010111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011010111100)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b10011010111101) && ({row_reg, col_reg}<14'b10011100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10011100000010) && ({row_reg, col_reg}<14'b10011100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011100000100) && ({row_reg, col_reg}<14'b10011100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011100000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011100001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011100001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011100001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10011100001110) && ({row_reg, col_reg}<14'b10011100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011100010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011100010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011100010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011100010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10011100010100) && ({row_reg, col_reg}<14'b10011100010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011100010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011100010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011100011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011100011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b10011100011101) && ({row_reg, col_reg}<14'b10011100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011100100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011100100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011100100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10011100100111) && ({row_reg, col_reg}<14'b10011100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011100101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011100101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011100101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011100101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011100110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10011100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011100110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011100110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b10011100110101) && ({row_reg, col_reg}<14'b10011100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011100111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10011100111011) && ({row_reg, col_reg}<14'b10011100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011101000001) && ({row_reg, col_reg}<14'b10011101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10011101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10011101001001) && ({row_reg, col_reg}<14'b10011101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011101001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011101001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10011101001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011101010010) && ({row_reg, col_reg}<14'b10011101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011101010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011101010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011101010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011101011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011101011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10011101011010) && ({row_reg, col_reg}<14'b10011101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011101100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10011101100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10011101100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011101100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011101100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10011101100101) && ({row_reg, col_reg}<14'b10011101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011101110010) && ({row_reg, col_reg}<14'b10011101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011101110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011101111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10011101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011101111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10011101111100) && ({row_reg, col_reg}<14'b10011101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011101111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011101111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10011110000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011110000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011110000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10011110000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011110000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10011110000111) && ({row_reg, col_reg}<14'b10011110010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10011110010010) && ({row_reg, col_reg}<14'b10011110010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10011110010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10011110010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011110010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10011110010111) && ({row_reg, col_reg}<14'b10011110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011110011100) && ({row_reg, col_reg}<14'b10011110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011110011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10011110100001) && ({row_reg, col_reg}<14'b10011110100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011110100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011110100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10011110100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011110100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011110101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10011110101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10011110101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10011110101100) && ({row_reg, col_reg}<14'b10011110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011110101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10011110110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011110110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10011110110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10011110110100) && ({row_reg, col_reg}<14'b10011110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10011110110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011110111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10011110111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10011110111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10011110111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10011110111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10011110111101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10011110111110) && ({row_reg, col_reg}<14'b10100000001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100000001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10100000001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10100000001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100000001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100000010001) && ({row_reg, col_reg}<14'b10100000010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100000011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10100000011010) && ({row_reg, col_reg}<14'b10100000011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100000011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10100000011101) && ({row_reg, col_reg}<14'b10100000011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100000100000) && ({row_reg, col_reg}<14'b10100000100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100000100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10100000100110) && ({row_reg, col_reg}<14'b10100000101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100000101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100000101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100000101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100000101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10100000110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10100000110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10100000110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100000110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=14'b10100000110101) && ({row_reg, col_reg}<14'b10100000110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10100000110111) && ({row_reg, col_reg}<14'b10100000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100000111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100000111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10100000111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100000111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100000111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100000111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b10100000111111) && ({row_reg, col_reg}<14'b10100001000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100001000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100001000010) && ({row_reg, col_reg}<14'b10100001000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100001000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10100001000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10100001000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100001001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100001001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100001001010) && ({row_reg, col_reg}<14'b10100001001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100001001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10100001001101) && ({row_reg, col_reg}<14'b10100001001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100001001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10100001010001) && ({row_reg, col_reg}<14'b10100001010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100001010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100001010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10100001010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100001010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100001011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10100001011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10100001011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=14'b10100001011011) && ({row_reg, col_reg}<14'b10100001011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100001011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100001011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10100001011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10100001100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100001100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10100001100101) && ({row_reg, col_reg}<14'b10100001111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100001111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10100001111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10100001111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100001111011) && ({row_reg, col_reg}<14'b10100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100001111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100001111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100001111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10100010000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10100010000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100010000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100010000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10100010000100) && ({row_reg, col_reg}<14'b10100010000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100010000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10100010000111) && ({row_reg, col_reg}<14'b10100010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100010100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100010100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10100010100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10100010101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10100010101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100010101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100010101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100010101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100010101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100010101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10100010101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10100010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100010110010) && ({row_reg, col_reg}<14'b10100010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100010111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100010111011) && ({row_reg, col_reg}<14'b10100010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100010111111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10100011000000) && ({row_reg, col_reg}<14'b10100100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100100001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100100001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10100100001101) && ({row_reg, col_reg}<14'b10100100001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10100100001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10100100010000) && ({row_reg, col_reg}<14'b10100100010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100100010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10100100010011) && ({row_reg, col_reg}<14'b10100100010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100100010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10100100010110) && ({row_reg, col_reg}<14'b10100100011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=14'b10100100011000) && ({row_reg, col_reg}<14'b10100100011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10100100011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100100011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100100011101) && ({row_reg, col_reg}<14'b10100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100100100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100100100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10100100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100100101001) && ({row_reg, col_reg}<14'b10100100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100100101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100100101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100100110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100100110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10100100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100100110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10100100110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b10100100110101) && ({row_reg, col_reg}<14'b10100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100100111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100100111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10100100111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10100100111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100100111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10100100111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b10100100111111) && ({row_reg, col_reg}<14'b10100101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100101000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10100101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10100101000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10100101001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100101001001) && ({row_reg, col_reg}<14'b10100101001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100101001110) && ({row_reg, col_reg}<14'b10100101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100101010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100101010010) && ({row_reg, col_reg}<14'b10100101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100101010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10100101010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100101011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100101011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10100101011011) && ({row_reg, col_reg}<14'b10100101011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10100101011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10100101011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100101011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100101100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10100101100001) && ({row_reg, col_reg}<14'b10100101100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10100101100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100101100101) && ({row_reg, col_reg}<14'b10100101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100101111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10100101111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100101111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100101111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10100101111101) && ({row_reg, col_reg}<14'b10100110000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100110000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=14'b10100110000011) && ({row_reg, col_reg}<14'b10100110000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10100110000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10100110000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100110000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100110001000) && ({row_reg, col_reg}<14'b10100110100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100110100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100110100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10100110100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10100110101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10100110101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10100110101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b10100110101011) && ({row_reg, col_reg}<14'b10100110101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10100110101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10100110101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10100110101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10100110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100110110001) && ({row_reg, col_reg}<14'b10100110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100110110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10100110111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10100110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10100110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10100110111011) && ({row_reg, col_reg}<14'b10100110111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10100110111111)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10100111000000) && ({row_reg, col_reg}<14'b10101000001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101000001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101000001001) && ({row_reg, col_reg}<14'b10101000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101000001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10101000001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10101000001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10101000001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=14'b10101000010000) && ({row_reg, col_reg}<14'b10101000011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10101000011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101000011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10101000011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10101000011011) && ({row_reg, col_reg}<14'b10101000100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10101000100000) && ({row_reg, col_reg}<14'b10101000100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101000100010) && ({row_reg, col_reg}<14'b10101000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101000100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101000100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10101000101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10101000101001) && ({row_reg, col_reg}<14'b10101000101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10101000101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10101000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10101000101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10101000101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101000101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10101000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101000110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10101000110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10101000110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10101000110100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b10101000110101) && ({row_reg, col_reg}<14'b10101000110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101000110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101000111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101000111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10101000111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10101000111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101000111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10101000111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b10101000111111) && ({row_reg, col_reg}<14'b10101001000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101001000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101001000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101001000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10101001000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101001001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101001001001) && ({row_reg, col_reg}<14'b10101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10101001010001) && ({row_reg, col_reg}<14'b10101001010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101001010011) && ({row_reg, col_reg}<14'b10101001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101001010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101001010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10101001011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10101001011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101001011010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101001011011) && ({row_reg, col_reg}<14'b10101001011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101001011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101001011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10101001100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10101001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10101001100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101001100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101001100100) && ({row_reg, col_reg}<14'b10101001111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101001111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10101001111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10101001111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10101001111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10101001111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10101001111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=14'b10101001111110) && ({row_reg, col_reg}<14'b10101010000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10101010000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10101010000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10101010000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10101010000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10101010000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101010000101) && ({row_reg, col_reg}<14'b10101010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101010101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10101010101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10101010101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10101010101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10101010101101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10101010101110) && ({row_reg, col_reg}<14'b10101100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101100001001) && ({row_reg, col_reg}<14'b10101100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101100011110) && ({row_reg, col_reg}<14'b10101100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101100100011) && ({row_reg, col_reg}<14'b10101100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101100100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10101100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101100101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101100101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==14'b10101100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==14'b10101100101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101100101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101100101110) && ({row_reg, col_reg}<14'b10101100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101100110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10101100110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10101100110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101100110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10101100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10101100110110) && ({row_reg, col_reg}<14'b10101100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101100111000) && ({row_reg, col_reg}<14'b10101100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10101100111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==14'b10101100111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101100111101) && ({row_reg, col_reg}<14'b10101100111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=14'b10101100111111) && ({row_reg, col_reg}<14'b10101101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10101101000001) && ({row_reg, col_reg}<14'b10101101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101101000011) && ({row_reg, col_reg}<14'b10101101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101101010000) && ({row_reg, col_reg}<14'b10101101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101101010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101101010100) && ({row_reg, col_reg}<14'b10101101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101101010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10101101011000) && ({row_reg, col_reg}<14'b10101101011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=14'b10101101011011) && ({row_reg, col_reg}<14'b10101101011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=14'b10101101011101) && ({row_reg, col_reg}<14'b10101101100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==14'b10101101100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10101101100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10101101100011) && ({row_reg, col_reg}<14'b10101101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101101111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10101101111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==14'b10101101111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101101111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==14'b10101101111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=14'b10101101111111) && ({row_reg, col_reg}<14'b10101110000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==14'b10101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==14'b10101110000010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10101110000011) && ({row_reg, col_reg}<14'b10101110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101110000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10101110001000) && ({row_reg, col_reg}<14'b10101110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10101110101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10101110101111)) color_data = 12'b001000100010;

		if(({row_reg, col_reg}>=14'b10101110110000) && ({row_reg, col_reg}<14'b10110000001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110000001011) && ({row_reg, col_reg}<14'b10110000001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110000001101) && ({row_reg, col_reg}<14'b10110000010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110000010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110000010011) && ({row_reg, col_reg}<14'b10110000010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10110000010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110000010110) && ({row_reg, col_reg}<14'b10110000011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110000011010) && ({row_reg, col_reg}<14'b10110000011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110000011101) && ({row_reg, col_reg}<14'b10110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110000101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110000101011) && ({row_reg, col_reg}<14'b10110000110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110000110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10110000110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110000110011) && ({row_reg, col_reg}<14'b10110000111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110000111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110000111001) && ({row_reg, col_reg}<14'b10110001000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110001000011) && ({row_reg, col_reg}<14'b10110001000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110001000101) && ({row_reg, col_reg}<14'b10110001000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110001000111) && ({row_reg, col_reg}<14'b10110001001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110001001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110001010000) && ({row_reg, col_reg}<14'b10110001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110001010011) && ({row_reg, col_reg}<14'b10110001010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110001010101) && ({row_reg, col_reg}<14'b10110001011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110001011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10110001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10110001011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b10110001011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==14'b10110001011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10110001011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10110001100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10110001100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110001100010) && ({row_reg, col_reg}<14'b10110010000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110010000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10110010000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110010000111) && ({row_reg, col_reg}<14'b10110010100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110010100110) && ({row_reg, col_reg}<14'b10110010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110010101010) && ({row_reg, col_reg}<14'b10110010101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10110010101101)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10110010101110) && ({row_reg, col_reg}<14'b10110100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110100001101) && ({row_reg, col_reg}<14'b10110100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110100001111) && ({row_reg, col_reg}<14'b10110100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110100011001) && ({row_reg, col_reg}<14'b10110100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110100011011) && ({row_reg, col_reg}<14'b10110100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110100011111) && ({row_reg, col_reg}<14'b10110100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110100100001) && ({row_reg, col_reg}<14'b10110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110100100101) && ({row_reg, col_reg}<14'b10110100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110100100111) && ({row_reg, col_reg}<14'b10110100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110100101101) && ({row_reg, col_reg}<14'b10110100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10110100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110100110000) && ({row_reg, col_reg}<14'b10110100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110100111001) && ({row_reg, col_reg}<14'b10110101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110101000010) && ({row_reg, col_reg}<14'b10110101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110101000100) && ({row_reg, col_reg}<14'b10110101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110101000110) && ({row_reg, col_reg}<14'b10110101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110101001000) && ({row_reg, col_reg}<14'b10110101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110101010001) && ({row_reg, col_reg}<14'b10110101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110101010101) && ({row_reg, col_reg}<14'b10110101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110101011000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==14'b10110101011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=14'b10110101011010) && ({row_reg, col_reg}<14'b10110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110101111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10110101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110101111100) && ({row_reg, col_reg}<14'b10110101111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10110101111110) && ({row_reg, col_reg}<14'b10110110000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10110110000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10110110000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110110000100) && ({row_reg, col_reg}<14'b10110110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10110110100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10110110100001) && ({row_reg, col_reg}<14'b10110110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10110110111010) && ({row_reg, col_reg}<14'b10110110111100)) color_data = 12'b000100010001;

		if(({row_reg, col_reg}>=14'b10110110111100) && ({row_reg, col_reg}<14'b10111000001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111000001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111000001010) && ({row_reg, col_reg}<14'b10111000011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111000011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111000011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111000100000) && ({row_reg, col_reg}<14'b10111000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111000100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111000100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111000101000) && ({row_reg, col_reg}<14'b10111000101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111000101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111000101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10111000101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111000101110) && ({row_reg, col_reg}<14'b10111000110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111000110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111000110001) && ({row_reg, col_reg}<14'b10111000110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111000110101) && ({row_reg, col_reg}<14'b10111000110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111000110111) && ({row_reg, col_reg}<14'b10111000111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111000111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111000111010) && ({row_reg, col_reg}<14'b10111000111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111000111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10111000111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111000111110) && ({row_reg, col_reg}<14'b10111001000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111001000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111001000011) && ({row_reg, col_reg}<14'b10111001001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111001001000) && ({row_reg, col_reg}<14'b10111001001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111001001010) && ({row_reg, col_reg}<14'b10111001001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111001001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111001001101) && ({row_reg, col_reg}<14'b10111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111001010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111001010001) && ({row_reg, col_reg}<14'b10111001010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111001010101) && ({row_reg, col_reg}<14'b10111001010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==14'b10111001010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111001011000) && ({row_reg, col_reg}<14'b10111001011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111001011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111001011101) && ({row_reg, col_reg}<14'b10111001100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111001100000) && ({row_reg, col_reg}<14'b10111001111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111001111100) && ({row_reg, col_reg}<14'b10111001111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111001111111) && ({row_reg, col_reg}<14'b10111010000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111010000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111010000011) && ({row_reg, col_reg}<14'b10111010000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111010000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10111010000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=14'b10111010001000) && ({row_reg, col_reg}<14'b10111010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111010101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10111010101111)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=14'b10111010110000) && ({row_reg, col_reg}<14'b10111100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111100001011) && ({row_reg, col_reg}<14'b10111100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111100001101) && ({row_reg, col_reg}<14'b10111100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111100001111) && ({row_reg, col_reg}<14'b10111100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b10111100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111100100100) && ({row_reg, col_reg}<14'b10111100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111100101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==14'b10111100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111100110001) && ({row_reg, col_reg}<14'b10111100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111100110100) && ({row_reg, col_reg}<14'b10111100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111100111010) && ({row_reg, col_reg}<14'b10111101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111101000100) && ({row_reg, col_reg}<14'b10111101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111101000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=14'b10111101001000) && ({row_reg, col_reg}<14'b10111101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111101011001) && ({row_reg, col_reg}<14'b10111101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111101100010) && ({row_reg, col_reg}<14'b10111101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111101100100) && ({row_reg, col_reg}<14'b10111101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=14'b10111101111001) && ({row_reg, col_reg}<14'b10111101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=14'b10111101111011) && ({row_reg, col_reg}<14'b10111110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b10111110000101)) color_data = 12'b000100010001;








		if(({row_reg, col_reg}>=14'b10111110000110) && ({row_reg, col_reg}<=14'b11011011000111)) color_data = 12'b000000000000;
	end
endmodule