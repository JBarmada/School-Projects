module title_rom
	(
		input wire clk,
		input wire [8:0] row,
		input wire [9:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [8:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=19'b0000000000000000000) && ({row_reg, col_reg}<19'b0000000001001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000000001001010000) && ({row_reg, col_reg}<19'b0000000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000000001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000000001001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000000010000000000) && ({row_reg, col_reg}<19'b0000000011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000000011001010000) && ({row_reg, col_reg}<19'b0000000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000000011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000000011001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000000100000000000) && ({row_reg, col_reg}<19'b0000000101001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000000101001010000) && ({row_reg, col_reg}<19'b0000000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000000101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000000101001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000000110000000000) && ({row_reg, col_reg}<19'b0000000111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000000111001010000) && ({row_reg, col_reg}<19'b0000000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000000111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000000111001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000001000000000000) && ({row_reg, col_reg}<19'b0000001001001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000001001001010000) && ({row_reg, col_reg}<19'b0000001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000001001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000001001001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000001010000000000) && ({row_reg, col_reg}<19'b0000001011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000001011001010000) && ({row_reg, col_reg}<19'b0000001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000001011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000001011001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000001100000000000) && ({row_reg, col_reg}<19'b0000001101001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000001101001010000) && ({row_reg, col_reg}<19'b0000001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000001101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000001101001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000001110000000000) && ({row_reg, col_reg}<19'b0000001111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000001111001010000) && ({row_reg, col_reg}<19'b0000001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000001111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000001111001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000010000000000000) && ({row_reg, col_reg}<19'b0000010001001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000010001001010000) && ({row_reg, col_reg}<19'b0000010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000010001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000010001001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000010010000000000) && ({row_reg, col_reg}<19'b0000010011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000010011001010000) && ({row_reg, col_reg}<19'b0000010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000010011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000010011001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000010100000000000) && ({row_reg, col_reg}<19'b0000010101001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000010101001010000) && ({row_reg, col_reg}<19'b0000010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000010101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000010101001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000010110000000000) && ({row_reg, col_reg}<19'b0000010111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000010111001010000) && ({row_reg, col_reg}<19'b0000010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000010111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000010111001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000011000000000000) && ({row_reg, col_reg}<19'b0000011001001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000011001001010000) && ({row_reg, col_reg}<19'b0000011001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000011001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000011001001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000011010000000000) && ({row_reg, col_reg}<19'b0000011011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000011011001010000) && ({row_reg, col_reg}<19'b0000011011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000011011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000011011001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000011100000000000) && ({row_reg, col_reg}<19'b0000011101001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000011101001010000) && ({row_reg, col_reg}<19'b0000011101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000011101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000011101001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000011110000000000) && ({row_reg, col_reg}<19'b0000011111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000011111001010000) && ({row_reg, col_reg}<19'b0000011111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000011111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000011111001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0000100000000000000) && ({row_reg, col_reg}<19'b0000100001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000100001001010001) && ({row_reg, col_reg}<19'b0000100001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000100001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000100001001010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0000100010000000000) && ({row_reg, col_reg}<19'b0000100010100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000100010100010001) && ({row_reg, col_reg}<19'b0000100010100011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0000100010100011111) && ({row_reg, col_reg}<19'b0000100011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000100011001010001) && ({row_reg, col_reg}<19'b0000100011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000100011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000100011001010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0000100100000000000) && ({row_reg, col_reg}<19'b0000100100100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000100100100010001) && ({row_reg, col_reg}<19'b0000100100100011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0000100100100011111) && ({row_reg, col_reg}<19'b0000100101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000100101001010001) && ({row_reg, col_reg}<19'b0000100101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000100101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000100101001010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0000100110000000000) && ({row_reg, col_reg}<19'b0000100110100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000100110100010001) && ({row_reg, col_reg}<19'b0000100110100011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0000100110100011111) && ({row_reg, col_reg}<19'b0000100111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000100111001010001) && ({row_reg, col_reg}<19'b0000100111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000100111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000100111001010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0000101000000000000) && ({row_reg, col_reg}<19'b0000101000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000101000100010001) && ({row_reg, col_reg}<19'b0000101000100011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0000101000100011111) && ({row_reg, col_reg}<19'b0000101001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000101001001010001) && ({row_reg, col_reg}<19'b0000101001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000101001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000101001001010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0000101010000000000) && ({row_reg, col_reg}<19'b0000101010100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000101010100010001) && ({row_reg, col_reg}<19'b0000101010100011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0000101010100011111) && ({row_reg, col_reg}<19'b0000101011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000101011001010001) && ({row_reg, col_reg}<19'b0000101011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000101011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000101011001010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0000101100000000000) && ({row_reg, col_reg}<19'b0000101100100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000101100100010001) && ({row_reg, col_reg}<19'b0000101100100011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0000101100100011111) && ({row_reg, col_reg}<19'b0000101101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000101101001010001) && ({row_reg, col_reg}<19'b0000101101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000101101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000101101001010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0000101110000000000) && ({row_reg, col_reg}<19'b0000101110100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000101110100010001) && ({row_reg, col_reg}<19'b0000101110100011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0000101110100011111) && ({row_reg, col_reg}<19'b0000101111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000101111001010001) && ({row_reg, col_reg}<19'b0000101111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000101111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b0000101111001010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0000110000000000000) && ({row_reg, col_reg}<19'b0000110000100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0000110000100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0000110000100001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110000100010000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==19'b0000110000100010001)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==19'b0000110000100010010)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==19'b0000110000100010011)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==19'b0000110000100010100)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0000110000100010101)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==19'b0000110000100010110)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==19'b0000110000100010111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==19'b0000110000100011000)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0000110000100011001)) color_data = 12'b110111001101;
		if(({row_reg, col_reg}==19'b0000110000100011010)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0000110000100011011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0000110000100011100)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0000110000100011101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0000110000100011110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000110000100011111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=19'b0000110000100100000) && ({row_reg, col_reg}<19'b0000110001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000110001001010001) && ({row_reg, col_reg}<19'b0000110001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000110001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0000110001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0000110010000000000) && ({row_reg, col_reg}<19'b0000110010100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0000110010100001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0000110010100001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110010100010000)) color_data = 12'b110111001101;
		if(({row_reg, col_reg}==19'b0000110010100010001)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0000110010100010010)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0000110010100010011)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==19'b0000110010100010100)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0000110010100010101)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0000110010100010110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==19'b0000110010100010111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==19'b0000110010100011000)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0000110010100011001)) color_data = 12'b110111001101;
		if(({row_reg, col_reg}==19'b0000110010100011010)) color_data = 12'b011101101000;
		if(({row_reg, col_reg}==19'b0000110010100011011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0000110010100011100)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0000110010100011101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0000110010100011110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000110010100011111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=19'b0000110010100100000) && ({row_reg, col_reg}<19'b0000110011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000110011001010001) && ({row_reg, col_reg}<19'b0000110011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000110011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0000110011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0000110100000000000) && ({row_reg, col_reg}<19'b0000110100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0000110100100001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0000110100100001111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==19'b0000110100100010000)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0000110100100010001)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==19'b0000110100100010010)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}==19'b0000110100100010011)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0000110100100010100)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==19'b0000110100100010101)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}>=19'b0000110100100010110) && ({row_reg, col_reg}<19'b0000110100100011000)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==19'b0000110100100011000)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0000110100100011001)) color_data = 12'b110110111101;
		if(({row_reg, col_reg}==19'b0000110100100011010)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==19'b0000110100100011011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0000110100100011100) && ({row_reg, col_reg}<19'b0000110100100011110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0000110100100011110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000110100100011111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=19'b0000110100100100000) && ({row_reg, col_reg}<19'b0000110101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000110101001010001) && ({row_reg, col_reg}<19'b0000110101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000110101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0000110101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0000110110000000000) && ({row_reg, col_reg}<19'b0000110110100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0000110110100001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0000110110100001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000110110100010000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==19'b0000110110100010001)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==19'b0000110110100010010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0000110110100010011)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==19'b0000110110100010100)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0000110110100010101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0000110110100010110) && ({row_reg, col_reg}<19'b0000110110100011000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000110110100011000)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0000110110100011001)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0000110110100011010)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}==19'b0000110110100011011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0000110110100011100) && ({row_reg, col_reg}<19'b0000110110100011110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0000110110100011110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000110110100011111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0000110110100100000) && ({row_reg, col_reg}<19'b0000110111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000110111001010001) && ({row_reg, col_reg}<19'b0000110111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000110111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0000110111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0000111000000000000) && ({row_reg, col_reg}<19'b0000111000100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0000111000100001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0000111000100001111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==19'b0000111000100010000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==19'b0000111000100010001)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=19'b0000111000100010010) && ({row_reg, col_reg}<19'b0000111000100010101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0000111000100010101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111000100010110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0000111000100010111)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0000111000100011000)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}==19'b0000111000100011001)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0000111000100011010)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==19'b0000111000100011011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111000100011100)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0000111000100011101)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0000111000100011110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111000100011111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0000111000100100000) && ({row_reg, col_reg}<19'b0000111001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000111001001010001) && ({row_reg, col_reg}<19'b0000111001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0000111001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0000111010000000000) && ({row_reg, col_reg}<19'b0000111010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0000111010100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0000111010100001100) && ({row_reg, col_reg}<19'b0000111010100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0000111010100001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0000111010100001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000111010100010000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==19'b0000111010100010001)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=19'b0000111010100010010) && ({row_reg, col_reg}<19'b0000111010100010100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0000111010100010100) && ({row_reg, col_reg}<19'b0000111010100010110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0000111010100010110)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0000111010100010111)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==19'b0000111010100011000)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}==19'b0000111010100011001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==19'b0000111010100011010)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}==19'b0000111010100011011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111010100011100)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0000111010100011101)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0000111010100011110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111010100011111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0000111010100100000) && ({row_reg, col_reg}<19'b0000111011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000111011001010001) && ({row_reg, col_reg}<19'b0000111011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0000111011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0000111100000000000) && ({row_reg, col_reg}<19'b0000111100100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0000111100100001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0000111100100001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0000111100100001100) && ({row_reg, col_reg}<19'b0000111100100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0000111100100001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0000111100100001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000111100100010000)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==19'b0000111100100010001)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0000111100100010010) && ({row_reg, col_reg}<19'b0000111100100010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111100100010110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0000111100100010111)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0000111100100011000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==19'b0000111100100011001)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0000111100100011010)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0000111100100011011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111100100011100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0000111100100011101)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==19'b0000111100100011110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111100100011111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0000111100100100000) && ({row_reg, col_reg}<19'b0000111101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000111101001010001) && ({row_reg, col_reg}<19'b0000111101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0000111101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0000111110000000000) && ({row_reg, col_reg}<19'b0000111110100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0000111110100001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0000111110100001001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==19'b0000111110100001010)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==19'b0000111110100001011)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==19'b0000111110100001100)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==19'b0000111110100001101)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==19'b0000111110100001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==19'b0000111110100001111)) color_data = 12'b110111001101;
		if(({row_reg, col_reg}==19'b0000111110100010000)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==19'b0000111110100010001)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0000111110100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0000111110100010011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0000111110100010100)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0000111110100010101) && ({row_reg, col_reg}<19'b0000111110100010111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0000111110100010111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0000111110100011000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==19'b0000111110100011001)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}==19'b0000111110100011010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==19'b0000111110100011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0000111110100011100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0000111110100011101)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=19'b0000111110100011110) && ({row_reg, col_reg}<19'b0000111110100100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0000111110100100000) && ({row_reg, col_reg}<19'b0000111111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0000111111001010001) && ({row_reg, col_reg}<19'b0000111111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0000111111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0000111111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001000000000000000) && ({row_reg, col_reg}<19'b0001000000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001000000100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001000000100000001) && ({row_reg, col_reg}<19'b0001000000100001000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001000000100001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001000000100001001)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==19'b0001000000100001010)) color_data = 12'b111010111100;
		if(({row_reg, col_reg}==19'b0001000000100001011)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}==19'b0001000000100001100)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}>=19'b0001000000100001101) && ({row_reg, col_reg}<19'b0001000000100001111)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==19'b0001000000100001111)) color_data = 12'b101001111000;
		if(({row_reg, col_reg}>=19'b0001000000100010000) && ({row_reg, col_reg}<19'b0001000000100010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001000000100010101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0001000000100010110)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==19'b0001000000100010111)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==19'b0001000000100011000)) color_data = 12'b110010011010;
		if(({row_reg, col_reg}==19'b0001000000100011001)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==19'b0001000000100011010)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0001000000100011011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001000000100011100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0001000000100011101) && ({row_reg, col_reg}<19'b0001000000100011111)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0001000000100011111)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0001000000100100000) && ({row_reg, col_reg}<19'b0001000001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001000001001010001) && ({row_reg, col_reg}<19'b0001000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001000001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001000001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001000010000000000) && ({row_reg, col_reg}<19'b0001000010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001000010100000000) && ({row_reg, col_reg}<19'b0001000010100001000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001000010100001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001000010100001001)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==19'b0001000010100001010)) color_data = 12'b110110101011;
		if(({row_reg, col_reg}==19'b0001000010100001011)) color_data = 12'b110010011010;
		if(({row_reg, col_reg}==19'b0001000010100001100)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==19'b0001000010100001101)) color_data = 12'b110010011010;
		if(({row_reg, col_reg}==19'b0001000010100001110)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==19'b0001000010100001111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==19'b0001000010100010000)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0001000010100010001)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==19'b0001000010100010010)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==19'b0001000010100010011)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==19'b0001000010100010100)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==19'b0001000010100010101)) color_data = 12'b100101100111;
		if(({row_reg, col_reg}==19'b0001000010100010110)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==19'b0001000010100010111)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==19'b0001000010100011000)) color_data = 12'b110110101011;
		if(({row_reg, col_reg}==19'b0001000010100011001)) color_data = 12'b100101100111;
		if(({row_reg, col_reg}==19'b0001000010100011010)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}>=19'b0001000010100011011) && ({row_reg, col_reg}<19'b0001000010100011101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0001000010100011101) && ({row_reg, col_reg}<19'b0001000010100011111)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0001000010100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001000010100100000) && ({row_reg, col_reg}<19'b0001000011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001000011001010001) && ({row_reg, col_reg}<19'b0001000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001000011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001000011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001000100000000000) && ({row_reg, col_reg}<19'b0001000100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001000100100000000) && ({row_reg, col_reg}<19'b0001000100100001000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001000100100001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001000100100001001)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==19'b0001000100100001010)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==19'b0001000100100001011)) color_data = 12'b110110101011;
		if(({row_reg, col_reg}>=19'b0001000100100001100) && ({row_reg, col_reg}<19'b0001000100100001110)) color_data = 12'b110010011010;
		if(({row_reg, col_reg}==19'b0001000100100001110)) color_data = 12'b100101100111;
		if(({row_reg, col_reg}==19'b0001000100100001111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==19'b0001000100100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001000100100010001)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==19'b0001000100100010010)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==19'b0001000100100010011)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}>=19'b0001000100100010100) && ({row_reg, col_reg}<19'b0001000100100010110)) color_data = 12'b110010011010;
		if(({row_reg, col_reg}==19'b0001000100100010110)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=19'b0001000100100010111) && ({row_reg, col_reg}<19'b0001000100100011001)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==19'b0001000100100011001)) color_data = 12'b100101100111;
		if(({row_reg, col_reg}==19'b0001000100100011010)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=19'b0001000100100011011) && ({row_reg, col_reg}<19'b0001000100100011101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0001000100100011101)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0001000100100011110)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001000100100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001000100100100000) && ({row_reg, col_reg}<19'b0001000101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001000101001010001) && ({row_reg, col_reg}<19'b0001000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001000101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001000101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001000110000000000) && ({row_reg, col_reg}<19'b0001000110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001000110100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001000110100000001) && ({row_reg, col_reg}<19'b0001000110100001000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001000110100001000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0001000110100001001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==19'b0001000110100001010)) color_data = 12'b110110111100;
		if(({row_reg, col_reg}==19'b0001000110100001011)) color_data = 12'b111010111100;
		if(({row_reg, col_reg}==19'b0001000110100001100)) color_data = 12'b110110101011;
		if(({row_reg, col_reg}==19'b0001000110100001101)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}==19'b0001000110100001110)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==19'b0001000110100001111)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==19'b0001000110100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001000110100010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==19'b0001000110100010010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==19'b0001000110100010011)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==19'b0001000110100010100)) color_data = 12'b111011001100;
		if(({row_reg, col_reg}==19'b0001000110100010101)) color_data = 12'b110110101011;
		if(({row_reg, col_reg}==19'b0001000110100010110)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==19'b0001000110100010111)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==19'b0001000110100011000)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==19'b0001000110100011001)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==19'b0001000110100011010)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}>=19'b0001000110100011011) && ({row_reg, col_reg}<19'b0001000110100011111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001000110100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001000110100100000) && ({row_reg, col_reg}<19'b0001000111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001000111001010001) && ({row_reg, col_reg}<19'b0001000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001000111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001000111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001001000000000000) && ({row_reg, col_reg}<19'b0001001000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001001000100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001001000100000001) && ({row_reg, col_reg}<19'b0001001000100001000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001001000100001000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0001001000100001001)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==19'b0001001000100001010)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==19'b0001001000100001011)) color_data = 12'b110010011010;
		if(({row_reg, col_reg}==19'b0001001000100001100)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==19'b0001001000100001101)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==19'b0001001000100001110)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=19'b0001001000100001111) && ({row_reg, col_reg}<19'b0001001000100010001)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0001001000100010001)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==19'b0001001000100010010)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}>=19'b0001001000100010011) && ({row_reg, col_reg}<19'b0001001000100010101)) color_data = 12'b111011001101;
		if(({row_reg, col_reg}==19'b0001001000100010101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==19'b0001001000100010110)) color_data = 12'b101001111000;
		if(({row_reg, col_reg}==19'b0001001000100010111)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==19'b0001001000100011000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==19'b0001001000100011001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0001001000100011010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0001001000100011011) && ({row_reg, col_reg}<19'b0001001000100011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001001000100011101) && ({row_reg, col_reg}<19'b0001001000100011111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001001000100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001001000100100000) && ({row_reg, col_reg}<19'b0001001001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001001001001010001) && ({row_reg, col_reg}<19'b0001001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001001001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001001001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001001010000000000) && ({row_reg, col_reg}<19'b0001001010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001001010100000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001001010100000001) && ({row_reg, col_reg}<19'b0001001010100001000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001001010100001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001001010100001001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0001001010100001010)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==19'b0001001010100001011)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==19'b0001001010100001100)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==19'b0001001010100001101)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==19'b0001001010100001110)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0001001010100001111) && ({row_reg, col_reg}<19'b0001001010100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001001010100010001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==19'b0001001010100010010)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==19'b0001001010100010011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==19'b0001001010100010100)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==19'b0001001010100010101)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==19'b0001001010100010110)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==19'b0001001010100010111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=19'b0001001010100011000) && ({row_reg, col_reg}<19'b0001001010100100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001001010100100000) && ({row_reg, col_reg}<19'b0001001011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001001011001010001) && ({row_reg, col_reg}<19'b0001001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001001011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001001011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001001100000000000) && ({row_reg, col_reg}<19'b0001001100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001001100100000000) && ({row_reg, col_reg}<19'b0001001100100001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001001100100001011) && ({row_reg, col_reg}<19'b0001001100100001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0001001100100001101) && ({row_reg, col_reg}<19'b0001001100100010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001001100100010010) && ({row_reg, col_reg}<19'b0001001100100010100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0001001100100010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0001001100100010101) && ({row_reg, col_reg}<19'b0001001100100100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001001100100100000) && ({row_reg, col_reg}<19'b0001001101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001001101001010001) && ({row_reg, col_reg}<19'b0001001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001001101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001001101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001001110000000000) && ({row_reg, col_reg}<19'b0001001110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001001110100000000) && ({row_reg, col_reg}<19'b0001001110100001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001001110100001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==19'b0001001110100001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001001110100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001001110100001011) && ({row_reg, col_reg}<19'b0001001110100010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001001110100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001001110100010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001001110100010010)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0001001110100010011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0001001110100010100) && ({row_reg, col_reg}<19'b0001001110100010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001001110100010110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0001001110100010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==19'b0001001110100011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001001110100011001)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0001001110100011010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==19'b0001001110100011011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0001001110100011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001001110100011101) && ({row_reg, col_reg}<19'b0001001111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001001111001010001) && ({row_reg, col_reg}<19'b0001001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001001111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001001111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001010000000000000) && ({row_reg, col_reg}<19'b0001010000101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001010000101110001) && ({row_reg, col_reg}<19'b0001010000101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001010000101110100) && ({row_reg, col_reg}<19'b0001010000110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001010000110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001010000110110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0001010000110110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0001010000110110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0001010000110110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001010000110110101) && ({row_reg, col_reg}<19'b0001010001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001010001001010001) && ({row_reg, col_reg}<19'b0001010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001010001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001010001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001010010000000000) && ({row_reg, col_reg}<19'b0001010010110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001010010110110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010010110110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010010110110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010010110110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010010110110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0001010010110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001010010110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001010010110110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001010010110111000) && ({row_reg, col_reg}<19'b0001010011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001010011001010001) && ({row_reg, col_reg}<19'b0001010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001010011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001010011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001010100000000000) && ({row_reg, col_reg}<19'b0001010100101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001010100101110011) && ({row_reg, col_reg}<19'b0001010100101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001010100101110110) && ({row_reg, col_reg}<19'b0001010100110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001010100110101110) && ({row_reg, col_reg}<19'b0001010100110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001010100110110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0001010100110110001) && ({row_reg, col_reg}<19'b0001010100110110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001010100110110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010100110110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0001010100110110101) && ({row_reg, col_reg}<19'b0001010101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001010101001010001) && ({row_reg, col_reg}<19'b0001010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001010101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001010101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001010110000000000) && ({row_reg, col_reg}<19'b0001010110101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001010110101110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001010110101110010) && ({row_reg, col_reg}<19'b0001010110101110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0001010110101110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0001010110101110101) && ({row_reg, col_reg}<19'b0001010110110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001010110110101110) && ({row_reg, col_reg}<19'b0001010110110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001010110110110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0001010110110110001) && ({row_reg, col_reg}<19'b0001010110110110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010110110110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010110110110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0001010110110110101) && ({row_reg, col_reg}<19'b0001010111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001010111001010001) && ({row_reg, col_reg}<19'b0001010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001010111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001010111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001011000000000000) && ({row_reg, col_reg}<19'b0001011000101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001011000101110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0001011000101110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011000101110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011000101110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0001011000101110101) && ({row_reg, col_reg}<19'b0001011000101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001011000101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001011000101111000) && ({row_reg, col_reg}<19'b0001011000110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001011000110101110) && ({row_reg, col_reg}<19'b0001011000110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001011000110110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011000110110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011000110110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011000110110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0001011000110110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001011000110110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001011000110110110) && ({row_reg, col_reg}<19'b0001011001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001011001001010001) && ({row_reg, col_reg}<19'b0001011001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001011001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001011001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001011010000000000) && ({row_reg, col_reg}<19'b0001011010101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001011010101110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0001011010101110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011010101110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011010101110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0001011010101110101) && ({row_reg, col_reg}<19'b0001011010110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001011010110101110) && ({row_reg, col_reg}<19'b0001011010110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001011010110110000) && ({row_reg, col_reg}<19'b0001011010110110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001011010110110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001011010110110100) && ({row_reg, col_reg}<19'b0001011011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001011011001010001) && ({row_reg, col_reg}<19'b0001011011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001011011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001011011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001011100000000000) && ({row_reg, col_reg}<19'b0001011100101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001011100101110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0001011100101110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011100101110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011100101110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011100101110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0001011100101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001011100101110111) && ({row_reg, col_reg}<19'b0001011101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001011101001010001) && ({row_reg, col_reg}<19'b0001011101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001011101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001011101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001011110000000000) && ({row_reg, col_reg}<19'b0001011110101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001011110101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0001011110101110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0001011110101110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0001011110101110011) && ({row_reg, col_reg}<19'b0001011110101110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001011110101110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011110101110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0001011110101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001011110101111000) && ({row_reg, col_reg}<19'b0001011110110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001011110110110000) && ({row_reg, col_reg}<19'b0001011110110110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001011110110110011) && ({row_reg, col_reg}<19'b0001011110110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001011110110110110) && ({row_reg, col_reg}<19'b0001011110110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001011110110111000) && ({row_reg, col_reg}<19'b0001011111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001011111001010001) && ({row_reg, col_reg}<19'b0001011111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001011111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001011111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001100000000000000) && ({row_reg, col_reg}<19'b0001100000010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100000010110001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001100000010110010) && ({row_reg, col_reg}<19'b0001100000010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100000010110111) && ({row_reg, col_reg}<19'b0001100000010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001100000010111001) && ({row_reg, col_reg}<19'b0001100000011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001100000011000000) && ({row_reg, col_reg}<19'b0001100000100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100000100100100) && ({row_reg, col_reg}<19'b0001100000100101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100000100101000)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0001100000100101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100000100101010) && ({row_reg, col_reg}<19'b0001100000101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100000101101010) && ({row_reg, col_reg}<19'b0001100000101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001100000101101100) && ({row_reg, col_reg}<19'b0001100000101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100000101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001100000101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100000101110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001100000101110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100000101110100) && ({row_reg, col_reg}<19'b0001100000101110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0001100000101110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0001100000101110111) && ({row_reg, col_reg}<19'b0001100000110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100000110001000) && ({row_reg, col_reg}<19'b0001100000110001010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0001100000110001010) && ({row_reg, col_reg}<19'b0001100000110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100000110001110) && ({row_reg, col_reg}<19'b0001100000110010000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0001100000110010000) && ({row_reg, col_reg}<19'b0001100001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100001001010001) && ({row_reg, col_reg}<19'b0001100001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001100001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001100010000000000) && ({row_reg, col_reg}<19'b0001100010010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100010010110000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100010010110001)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}==19'b0001100010010110010)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0001100010010110011)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0001100010010110100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100010010110101) && ({row_reg, col_reg}<19'b0001100010010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100010010110111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0001100010010111000) && ({row_reg, col_reg}<19'b0001100010011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001100010011000000) && ({row_reg, col_reg}<19'b0001100010100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100010100100100) && ({row_reg, col_reg}<19'b0001100010100100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100010100100110) && ({row_reg, col_reg}<19'b0001100010100101000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001100010100101000)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}>=19'b0001100010100101001) && ({row_reg, col_reg}<19'b0001100010100101011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100010100101011) && ({row_reg, col_reg}<19'b0001100010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100010100101110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0001100010100101111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0001100010100110000) && ({row_reg, col_reg}<19'b0001100010101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100010101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0001100010101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100010101110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100010101110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0001100010101110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0001100010101110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001100010101110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001100010101110111) && ({row_reg, col_reg}<19'b0001100010110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100010110001000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100010110001001) && ({row_reg, col_reg}<19'b0001100010110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100010110001110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100010110001111)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0001100010110010000) && ({row_reg, col_reg}<19'b0001100011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100011001010001) && ({row_reg, col_reg}<19'b0001100011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001100011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001100100000000000) && ({row_reg, col_reg}<19'b0001100100010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100100010110000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100100010110001)) color_data = 12'b000100100100;
		if(({row_reg, col_reg}>=19'b0001100100010110010) && ({row_reg, col_reg}<19'b0001100100010110100)) color_data = 12'b001101000110;
		if(({row_reg, col_reg}==19'b0001100100010110100)) color_data = 12'b001000110101;
		if(({row_reg, col_reg}==19'b0001100100010110101)) color_data = 12'b000100010011;
		if(({row_reg, col_reg}==19'b0001100100010110110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100100010110111) && ({row_reg, col_reg}<19'b0001100100010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100100010111100) && ({row_reg, col_reg}<19'b0001100100011000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001100100011000000) && ({row_reg, col_reg}<19'b0001100100100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100100100100100) && ({row_reg, col_reg}<19'b0001100100100100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100100100100110) && ({row_reg, col_reg}<19'b0001100100100101010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001100100100101010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100100100101011) && ({row_reg, col_reg}<19'b0001100100100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100100100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0001100100100101111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=19'b0001100100100110000) && ({row_reg, col_reg}<19'b0001100100101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100100101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001100100101101001) && ({row_reg, col_reg}<19'b0001100100101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100100101110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0001100100101110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100100101110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100100101110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0001100100101110100) && ({row_reg, col_reg}<19'b0001100100101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100100101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001100100101110111) && ({row_reg, col_reg}<19'b0001100101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100101001010001) && ({row_reg, col_reg}<19'b0001100101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001100101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001100110000000000) && ({row_reg, col_reg}<19'b0001100110010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100110010101111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100110010110000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001100110010110001)) color_data = 12'b000000100101;
		if(({row_reg, col_reg}==19'b0001100110010110010)) color_data = 12'b001101011000;
		if(({row_reg, col_reg}==19'b0001100110010110011)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==19'b0001100110010110100)) color_data = 12'b010001011000;
		if(({row_reg, col_reg}==19'b0001100110010110101)) color_data = 12'b001000110101;
		if(({row_reg, col_reg}==19'b0001100110010110110)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0001100110010110111) && ({row_reg, col_reg}<19'b0001100110010111001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100110010111001) && ({row_reg, col_reg}<19'b0001100110100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100110100100100) && ({row_reg, col_reg}<19'b0001100110100100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001100110100100110) && ({row_reg, col_reg}<19'b0001100110100101000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001100110100101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100110100101001)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0001100110100101010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0001100110100101011) && ({row_reg, col_reg}<19'b0001100110100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100110100101110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0001100110100101111)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}>=19'b0001100110100110000) && ({row_reg, col_reg}<19'b0001100110101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100110101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001100110101101001) && ({row_reg, col_reg}<19'b0001100110101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001100110101101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001100110101101110) && ({row_reg, col_reg}<19'b0001100110101110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001100110101110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100110101110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100110101110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0001100110101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001100110101110100) && ({row_reg, col_reg}<19'b0001100111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001100111001010001) && ({row_reg, col_reg}<19'b0001100111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001100111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001100111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001101000000000000) && ({row_reg, col_reg}<19'b0001101000010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101000010101111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001101000010110000)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0001101000010110001)) color_data = 12'b000000010111;
		if(({row_reg, col_reg}==19'b0001101000010110010)) color_data = 12'b001001011010;
		if(({row_reg, col_reg}==19'b0001101000010110011)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==19'b0001101000010110100)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==19'b0001101000010110101)) color_data = 12'b001000110111;
		if(({row_reg, col_reg}==19'b0001101000010110110)) color_data = 12'b000000010100;
		if(({row_reg, col_reg}>=19'b0001101000010110111) && ({row_reg, col_reg}<19'b0001101000010111001)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001101000010111001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001101000010111010) && ({row_reg, col_reg}<19'b0001101000100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001101000100100100) && ({row_reg, col_reg}<19'b0001101000100100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001101000100100110) && ({row_reg, col_reg}<19'b0001101000100101000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001101000100101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001101000100101001)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0001101000100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001101000100101011) && ({row_reg, col_reg}<19'b0001101000100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101000100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0001101000100101110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0001101000100101111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001101000100110000) && ({row_reg, col_reg}<19'b0001101000101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101000101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001101000101101001) && ({row_reg, col_reg}<19'b0001101000101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101000101101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001101000101101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0001101000101101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101000101101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101000101110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101000101110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101000101110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0001101000101110011) && ({row_reg, col_reg}<19'b0001101001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001101001001010001) && ({row_reg, col_reg}<19'b0001101001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001101001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001101001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001101010000000000) && ({row_reg, col_reg}<19'b0001101010010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101010010101111)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001101010010110000)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==19'b0001101010010110001)) color_data = 12'b000000011000;
		if(({row_reg, col_reg}==19'b0001101010010110010)) color_data = 12'b001001001011;
		if(({row_reg, col_reg}==19'b0001101010010110011)) color_data = 12'b010001101101;
		if(({row_reg, col_reg}==19'b0001101010010110100)) color_data = 12'b001101101100;
		if(({row_reg, col_reg}==19'b0001101010010110101)) color_data = 12'b001001001001;
		if(({row_reg, col_reg}==19'b0001101010010110110)) color_data = 12'b000000110111;
		if(({row_reg, col_reg}==19'b0001101010010110111)) color_data = 12'b000000100101;
		if(({row_reg, col_reg}==19'b0001101010010111000)) color_data = 12'b000000010100;
		if(({row_reg, col_reg}==19'b0001101010010111001)) color_data = 12'b000000010011;
		if(({row_reg, col_reg}==19'b0001101010010111010)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}==19'b0001101010010111011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0001101010010111100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001101010010111101) && ({row_reg, col_reg}<19'b0001101010100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001101010100100100) && ({row_reg, col_reg}<19'b0001101010100101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001101010100101001)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0001101010100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001101010100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101010100101100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0001101010100101101)) color_data = 12'b010101010010;
		if(({row_reg, col_reg}==19'b0001101010100101110)) color_data = 12'b010101100001;
		if(({row_reg, col_reg}==19'b0001101010100101111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=19'b0001101010100110000) && ({row_reg, col_reg}<19'b0001101010101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101010101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0001101010101101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0001101010101101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0001101010101101110) && ({row_reg, col_reg}<19'b0001101010101110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101010101110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101010101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101010101110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0001101010101110011) && ({row_reg, col_reg}<19'b0001101010110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101010110001010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0001101010110001011) && ({row_reg, col_reg}<19'b0001101010110001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==19'b0001101010110001101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001101010110001110) && ({row_reg, col_reg}<19'b0001101011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001101011001010001) && ({row_reg, col_reg}<19'b0001101011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001101011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001101011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001101100000000000) && ({row_reg, col_reg}<19'b0001101100010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101100010101111)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001101100010110000)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==19'b0001101100010110001)) color_data = 12'b000000101011;
		if(({row_reg, col_reg}==19'b0001101100010110010)) color_data = 12'b000101001101;
		if(({row_reg, col_reg}==19'b0001101100010110011)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==19'b0001101100010110100)) color_data = 12'b001101101101;
		if(({row_reg, col_reg}==19'b0001101100010110101)) color_data = 12'b001101011100;
		if(({row_reg, col_reg}==19'b0001101100010110110)) color_data = 12'b001101011011;
		if(({row_reg, col_reg}==19'b0001101100010110111)) color_data = 12'b001101011010;
		if(({row_reg, col_reg}==19'b0001101100010111000)) color_data = 12'b000000110110;
		if(({row_reg, col_reg}==19'b0001101100010111001)) color_data = 12'b000000110101;
		if(({row_reg, col_reg}==19'b0001101100010111010)) color_data = 12'b000000100011;
		if(({row_reg, col_reg}==19'b0001101100010111011)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}==19'b0001101100010111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0001101100010111101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001101100010111110) && ({row_reg, col_reg}<19'b0001101100100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001101100100100100) && ({row_reg, col_reg}<19'b0001101100100101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001101100100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001101100100101010) && ({row_reg, col_reg}<19'b0001101100100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101100100101100)) color_data = 12'b010001000001;
		if(({row_reg, col_reg}==19'b0001101100100101101)) color_data = 12'b101010110111;
		if(({row_reg, col_reg}==19'b0001101100100101110)) color_data = 12'b101010110110;
		if(({row_reg, col_reg}==19'b0001101100100101111)) color_data = 12'b010101100010;
		if(({row_reg, col_reg}>=19'b0001101100100110000) && ({row_reg, col_reg}<19'b0001101100101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101100101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001101100101101001) && ({row_reg, col_reg}<19'b0001101100101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101100101101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001101100101101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101100101101101) && ({row_reg, col_reg}<19'b0001101100101101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101100101101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101100101110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101100101110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0001101100101110010) && ({row_reg, col_reg}<19'b0001101100110001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101100110001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001101100110001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0001101100110001011) && ({row_reg, col_reg}<19'b0001101100110001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==19'b0001101100110001101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==19'b0001101100110001110)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001101100110001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001101100110010000) && ({row_reg, col_reg}<19'b0001101101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001101101001010001) && ({row_reg, col_reg}<19'b0001101101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001101101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001101101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001101110000000000) && ({row_reg, col_reg}<19'b0001101110010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101110010101111)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001101110010110000)) color_data = 12'b000000011000;
		if(({row_reg, col_reg}==19'b0001101110010110001)) color_data = 12'b000000101100;
		if(({row_reg, col_reg}==19'b0001101110010110010)) color_data = 12'b000101001110;
		if(({row_reg, col_reg}==19'b0001101110010110011)) color_data = 12'b001101011111;
		if(({row_reg, col_reg}==19'b0001101110010110100)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==19'b0001101110010110101)) color_data = 12'b001101101101;
		if(({row_reg, col_reg}==19'b0001101110010110110)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==19'b0001101110010110111)) color_data = 12'b010110001101;
		if(({row_reg, col_reg}==19'b0001101110010111000)) color_data = 12'b000101000111;
		if(({row_reg, col_reg}==19'b0001101110010111001)) color_data = 12'b000100110110;
		if(({row_reg, col_reg}==19'b0001101110010111010)) color_data = 12'b000100110100;
		if(({row_reg, col_reg}==19'b0001101110010111011)) color_data = 12'b000000100011;
		if(({row_reg, col_reg}==19'b0001101110010111100)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0001101110010111101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001101110010111110) && ({row_reg, col_reg}<19'b0001101110100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001101110100100100) && ({row_reg, col_reg}<19'b0001101110100101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001101110100101000) && ({row_reg, col_reg}<19'b0001101110100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101110100101100)) color_data = 12'b011001110011;
		if(({row_reg, col_reg}==19'b0001101110100101101)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==19'b0001101110100101110)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}==19'b0001101110100101111)) color_data = 12'b100010010100;
		if(({row_reg, col_reg}>=19'b0001101110100110000) && ({row_reg, col_reg}<19'b0001101110101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101110101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001101110101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101110101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001101110101101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0001101110101101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101110101101101) && ({row_reg, col_reg}<19'b0001101110101101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101110101101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101110101110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101110101110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0001101110101110010) && ({row_reg, col_reg}<19'b0001101110110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001101110110001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001101110110001001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==19'b0001101110110001010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=19'b0001101110110001011) && ({row_reg, col_reg}<19'b0001101110110001101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==19'b0001101110110001101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==19'b0001101110110001110)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001101110110001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001101110110010000) && ({row_reg, col_reg}<19'b0001101111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001101111001010001) && ({row_reg, col_reg}<19'b0001101111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001101111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001101111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001110000000000000) && ({row_reg, col_reg}<19'b0001110000010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110000010101010) && ({row_reg, col_reg}<19'b0001110000010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001110000010101100) && ({row_reg, col_reg}<19'b0001110000010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110000010101111)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001110000010110000)) color_data = 12'b000000011001;
		if(({row_reg, col_reg}==19'b0001110000010110001)) color_data = 12'b000000111110;
		if(({row_reg, col_reg}==19'b0001110000010110010)) color_data = 12'b001101011111;
		if(({row_reg, col_reg}>=19'b0001110000010110011) && ({row_reg, col_reg}<19'b0001110000010110101)) color_data = 12'b001001011110;
		if(({row_reg, col_reg}==19'b0001110000010110101)) color_data = 12'b010001111110;
		if(({row_reg, col_reg}==19'b0001110000010110110)) color_data = 12'b010001101101;
		if(({row_reg, col_reg}==19'b0001110000010110111)) color_data = 12'b001001011010;
		if(({row_reg, col_reg}==19'b0001110000010111000)) color_data = 12'b010110001100;
		if(({row_reg, col_reg}==19'b0001110000010111001)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==19'b0001110000010111010)) color_data = 12'b001101010110;
		if(({row_reg, col_reg}==19'b0001110000010111011)) color_data = 12'b000100110100;
		if(({row_reg, col_reg}==19'b0001110000010111100)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}==19'b0001110000010111101)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0001110000010111110) && ({row_reg, col_reg}<19'b0001110000011000000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001110000011000000) && ({row_reg, col_reg}<19'b0001110000011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110000011110110) && ({row_reg, col_reg}<19'b0001110000011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001110000011111000) && ({row_reg, col_reg}<19'b0001110000100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110000100100011) && ({row_reg, col_reg}<19'b0001110000100101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001110000100101000)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0001110000100101001) && ({row_reg, col_reg}<19'b0001110000100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110000100101011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0001110000100101100)) color_data = 12'b011101110011;
		if(({row_reg, col_reg}==19'b0001110000100101101)) color_data = 12'b110111101000;
		if(({row_reg, col_reg}==19'b0001110000100101110)) color_data = 12'b110111100111;
		if(({row_reg, col_reg}==19'b0001110000100101111)) color_data = 12'b100110100101;
		if(({row_reg, col_reg}>=19'b0001110000100110000) && ({row_reg, col_reg}<19'b0001110000101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110000101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0001110000101101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0001110000101101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001110000101101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001110000101101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110000101110000) && ({row_reg, col_reg}<19'b0001110000110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110000110000111) && ({row_reg, col_reg}<19'b0001110000110001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001110000110001010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001110000110001011)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==19'b0001110000110001100)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==19'b0001110000110001101)) color_data = 12'b011101000100;
		if(({row_reg, col_reg}==19'b0001110000110001110)) color_data = 12'b010000010001;
		if(({row_reg, col_reg}>=19'b0001110000110001111) && ({row_reg, col_reg}<19'b0001110000110010001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001110000110010001) && ({row_reg, col_reg}<19'b0001110000110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001110000110010101) && ({row_reg, col_reg}<19'b0001110001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110001001010001) && ({row_reg, col_reg}<19'b0001110001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001110001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001110001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001110010000000000) && ({row_reg, col_reg}<19'b0001110010010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110010010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001110010010101111)) color_data = 12'b000100010100;
		if(({row_reg, col_reg}==19'b0001110010010110000)) color_data = 12'b000100111011;
		if(({row_reg, col_reg}==19'b0001110010010110001)) color_data = 12'b001101101111;
		if(({row_reg, col_reg}==19'b0001110010010110010)) color_data = 12'b010001111111;
		if(({row_reg, col_reg}==19'b0001110010010110011)) color_data = 12'b001101101111;
		if(({row_reg, col_reg}==19'b0001110010010110100)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==19'b0001110010010110101)) color_data = 12'b010001111110;
		if(({row_reg, col_reg}==19'b0001110010010110110)) color_data = 12'b010001101101;
		if(({row_reg, col_reg}==19'b0001110010010110111)) color_data = 12'b001001011010;
		if(({row_reg, col_reg}==19'b0001110010010111000)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==19'b0001110010010111001)) color_data = 12'b001101011000;
		if(({row_reg, col_reg}==19'b0001110010010111010)) color_data = 12'b000100110101;
		if(({row_reg, col_reg}==19'b0001110010010111011)) color_data = 12'b000000100011;
		if(({row_reg, col_reg}==19'b0001110010010111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0001110010010111101) && ({row_reg, col_reg}<19'b0001110010010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110010010111111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001110010011000000) && ({row_reg, col_reg}<19'b0001110010100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110010100100011) && ({row_reg, col_reg}<19'b0001110010100100111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001110010100100111) && ({row_reg, col_reg}<19'b0001110010100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110010100101011)) color_data = 12'b001100110000;
		if(({row_reg, col_reg}==19'b0001110010100101100)) color_data = 12'b100110100101;
		if(({row_reg, col_reg}==19'b0001110010100101101)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==19'b0001110010100101110)) color_data = 12'b111011110111;
		if(({row_reg, col_reg}==19'b0001110010100101111)) color_data = 12'b100110100100;
		if(({row_reg, col_reg}==19'b0001110010100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110010100110001) && ({row_reg, col_reg}<19'b0001110010100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001110010100110100) && ({row_reg, col_reg}<19'b0001110010101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110010101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001110010101101001) && ({row_reg, col_reg}<19'b0001110010101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110010101101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001110010101101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0001110010101101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001110010101101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001110010101110000) && ({row_reg, col_reg}<19'b0001110010110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110010110000111) && ({row_reg, col_reg}<19'b0001110010110001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001110010110001010)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0001110010110001011)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}==19'b0001110010110001100)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==19'b0001110010110001101)) color_data = 12'b100001000100;
		if(({row_reg, col_reg}==19'b0001110010110001110)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==19'b0001110010110001111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001110010110010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001110010110010001) && ({row_reg, col_reg}<19'b0001110011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110011001010001) && ({row_reg, col_reg}<19'b0001110011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001110011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001110011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001110100000000000) && ({row_reg, col_reg}<19'b0001110100010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110100010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001110100010101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001110100010101111)) color_data = 12'b010001000110;
		if(({row_reg, col_reg}==19'b0001110100010110000)) color_data = 12'b010001101101;
		if(({row_reg, col_reg}==19'b0001110100010110001)) color_data = 12'b010101111111;
		if(({row_reg, col_reg}==19'b0001110100010110010)) color_data = 12'b011010001111;
		if(({row_reg, col_reg}==19'b0001110100010110011)) color_data = 12'b010101111111;
		if(({row_reg, col_reg}==19'b0001110100010110100)) color_data = 12'b010001101110;
		if(({row_reg, col_reg}==19'b0001110100010110101)) color_data = 12'b010101111110;
		if(({row_reg, col_reg}==19'b0001110100010110110)) color_data = 12'b010101101101;
		if(({row_reg, col_reg}==19'b0001110100010110111)) color_data = 12'b001101001001;
		if(({row_reg, col_reg}==19'b0001110100010111000)) color_data = 12'b000100110111;
		if(({row_reg, col_reg}==19'b0001110100010111001)) color_data = 12'b000100100101;
		if(({row_reg, col_reg}==19'b0001110100010111010)) color_data = 12'b000000010100;
		if(({row_reg, col_reg}==19'b0001110100010111011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001110100010111100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001110100010111101) && ({row_reg, col_reg}<19'b0001110100100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110100100100011) && ({row_reg, col_reg}<19'b0001110100100100111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001110100100100111) && ({row_reg, col_reg}<19'b0001110100100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110100100101001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0001110100100101010)) color_data = 12'b001101000001;
		if(({row_reg, col_reg}==19'b0001110100100101011)) color_data = 12'b011110000011;
		if(({row_reg, col_reg}==19'b0001110100100101100)) color_data = 12'b110111100111;
		if(({row_reg, col_reg}==19'b0001110100100101101)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==19'b0001110100100101110)) color_data = 12'b111011110111;
		if(({row_reg, col_reg}==19'b0001110100100101111)) color_data = 12'b101010110101;
		if(({row_reg, col_reg}==19'b0001110100100110000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001110100100110001) && ({row_reg, col_reg}<19'b0001110100101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110100101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001110100101101001) && ({row_reg, col_reg}<19'b0001110100101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110100101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001110100101101110) && ({row_reg, col_reg}<19'b0001110100110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110100110000000) && ({row_reg, col_reg}<19'b0001110100110000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001110100110000011) && ({row_reg, col_reg}<19'b0001110100110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110100110000111) && ({row_reg, col_reg}<19'b0001110100110001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001110100110001001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001110100110001010)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==19'b0001110100110001011)) color_data = 12'b011100110010;
		if(({row_reg, col_reg}==19'b0001110100110001100)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}==19'b0001110100110001101)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==19'b0001110100110001110)) color_data = 12'b010100000000;
		if(({row_reg, col_reg}==19'b0001110100110001111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0001110100110010000) && ({row_reg, col_reg}<19'b0001110101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110101001010001) && ({row_reg, col_reg}<19'b0001110101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001110101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001110101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001110110000000000) && ({row_reg, col_reg}<19'b0001110110010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110110010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001110110010101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001110110010101111)) color_data = 12'b010101010111;
		if(({row_reg, col_reg}==19'b0001110110010110000)) color_data = 12'b010001011011;
		if(({row_reg, col_reg}>=19'b0001110110010110001) && ({row_reg, col_reg}<19'b0001110110010110011)) color_data = 12'b010101111110;
		if(({row_reg, col_reg}==19'b0001110110010110011)) color_data = 12'b010001101101;
		if(({row_reg, col_reg}==19'b0001110110010110100)) color_data = 12'b010101101101;
		if(({row_reg, col_reg}==19'b0001110110010110101)) color_data = 12'b011001111110;
		if(({row_reg, col_reg}==19'b0001110110010110110)) color_data = 12'b010101111100;
		if(({row_reg, col_reg}==19'b0001110110010110111)) color_data = 12'b001101001001;
		if(({row_reg, col_reg}==19'b0001110110010111000)) color_data = 12'b000000010101;
		if(({row_reg, col_reg}==19'b0001110110010111001)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0001110110010111010)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0001110110010111011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0001110110010111100) && ({row_reg, col_reg}<19'b0001110110011000000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001110110011000000) && ({row_reg, col_reg}<19'b0001110110100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110110100100010) && ({row_reg, col_reg}<19'b0001110110100100111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001110110100100111) && ({row_reg, col_reg}<19'b0001110110100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110110100101001)) color_data = 12'b001101000010;
		if(({row_reg, col_reg}==19'b0001110110100101010)) color_data = 12'b100110100110;
		if(({row_reg, col_reg}==19'b0001110110100101011)) color_data = 12'b110111011000;
		if(({row_reg, col_reg}==19'b0001110110100101100)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}==19'b0001110110100101101)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==19'b0001110110100101110)) color_data = 12'b111011110111;
		if(({row_reg, col_reg}==19'b0001110110100101111)) color_data = 12'b110011010110;
		if(({row_reg, col_reg}==19'b0001110110100110000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==19'b0001110110100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001110110100110010) && ({row_reg, col_reg}<19'b0001110110100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110110100110110) && ({row_reg, col_reg}<19'b0001110110100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001110110100111000) && ({row_reg, col_reg}<19'b0001110110101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001110110101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001110110101101001) && ({row_reg, col_reg}<19'b0001110110101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110110101101100) && ({row_reg, col_reg}<19'b0001110110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001110110101101110) && ({row_reg, col_reg}<19'b0001110110110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110110110000000) && ({row_reg, col_reg}<19'b0001110110110000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001110110110000011) && ({row_reg, col_reg}<19'b0001110110110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110110110000110) && ({row_reg, col_reg}<19'b0001110110110001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001110110110001000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001110110110001001)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0001110110110001010)) color_data = 12'b010100100001;
		if(({row_reg, col_reg}==19'b0001110110110001011)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==19'b0001110110110001100)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}==19'b0001110110110001101)) color_data = 12'b100000110011;
		if(({row_reg, col_reg}==19'b0001110110110001110)) color_data = 12'b010100000000;
		if(({row_reg, col_reg}==19'b0001110110110001111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0001110110110010000) && ({row_reg, col_reg}<19'b0001110111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001110111001010001) && ({row_reg, col_reg}<19'b0001110111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001110111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001110111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001111000000000000) && ({row_reg, col_reg}<19'b0001111000010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111000010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111000010101010) && ({row_reg, col_reg}<19'b0001111000010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111000010101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0001111000010101111)) color_data = 12'b001101000101;
		if(({row_reg, col_reg}==19'b0001111000010110000)) color_data = 12'b001000110111;
		if(({row_reg, col_reg}==19'b0001111000010110001)) color_data = 12'b001001001010;
		if(({row_reg, col_reg}==19'b0001111000010110010)) color_data = 12'b001000111010;
		if(({row_reg, col_reg}==19'b0001111000010110011)) color_data = 12'b001000111001;
		if(({row_reg, col_reg}==19'b0001111000010110100)) color_data = 12'b010001011010;
		if(({row_reg, col_reg}==19'b0001111000010110101)) color_data = 12'b011101111100;
		if(({row_reg, col_reg}==19'b0001111000010110110)) color_data = 12'b011001111011;
		if(({row_reg, col_reg}==19'b0001111000010110111)) color_data = 12'b010001001000;
		if(({row_reg, col_reg}==19'b0001111000010111000)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}>=19'b0001111000010111001) && ({row_reg, col_reg}<19'b0001111000010111011)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}>=19'b0001111000010111011) && ({row_reg, col_reg}<19'b0001111000010111101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0001111000010111101) && ({row_reg, col_reg}<19'b0001111000011000000)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0001111000011000000) && ({row_reg, col_reg}<19'b0001111000100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111000100100010) && ({row_reg, col_reg}<19'b0001111000100100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001111000100100110) && ({row_reg, col_reg}<19'b0001111000100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111000100101001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==19'b0001111000100101010)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==19'b0001111000100101011)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0001111000100101100)) color_data = 12'b111011111000;
		if(({row_reg, col_reg}==19'b0001111000100101101)) color_data = 12'b110111110110;
		if(({row_reg, col_reg}==19'b0001111000100101110)) color_data = 12'b111011110110;
		if(({row_reg, col_reg}==19'b0001111000100101111)) color_data = 12'b111011111000;
		if(({row_reg, col_reg}==19'b0001111000100110000)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==19'b0001111000100110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111000100110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0001111000100110011) && ({row_reg, col_reg}<19'b0001111000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111000100110110) && ({row_reg, col_reg}<19'b0001111000100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111000100111000) && ({row_reg, col_reg}<19'b0001111000101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111000101101100) && ({row_reg, col_reg}<19'b0001111000101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111000101110000) && ({row_reg, col_reg}<19'b0001111000110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111000110000000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0001111000110000001) && ({row_reg, col_reg}<19'b0001111000110000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001111000110000011) && ({row_reg, col_reg}<19'b0001111000110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111000110000110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0001111000110000111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0001111000110001000)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==19'b0001111000110001001)) color_data = 12'b010100010000;
		if(({row_reg, col_reg}==19'b0001111000110001010)) color_data = 12'b011100110010;
		if(({row_reg, col_reg}==19'b0001111000110001011)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==19'b0001111000110001100)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==19'b0001111000110001101)) color_data = 12'b100000110010;
		if(({row_reg, col_reg}==19'b0001111000110001110)) color_data = 12'b011000010000;
		if(({row_reg, col_reg}==19'b0001111000110001111)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0001111000110010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001111000110010001) && ({row_reg, col_reg}<19'b0001111001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111001001010001) && ({row_reg, col_reg}<19'b0001111001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001111001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001111001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001111010000000000) && ({row_reg, col_reg}<19'b0001111010010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111010010101001) && ({row_reg, col_reg}<19'b0001111010010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111010010101011) && ({row_reg, col_reg}<19'b0001111010010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111010010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001111010010101111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==19'b0001111010010110000)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0001111010010110001)) color_data = 12'b000000010101;
		if(({row_reg, col_reg}>=19'b0001111010010110010) && ({row_reg, col_reg}<19'b0001111010010110100)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==19'b0001111010010110100)) color_data = 12'b001100111000;
		if(({row_reg, col_reg}==19'b0001111010010110101)) color_data = 12'b011001101011;
		if(({row_reg, col_reg}==19'b0001111010010110110)) color_data = 12'b011001101010;
		if(({row_reg, col_reg}==19'b0001111010010110111)) color_data = 12'b010001001000;
		if(({row_reg, col_reg}==19'b0001111010010111000)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}>=19'b0001111010010111001) && ({row_reg, col_reg}<19'b0001111010010111101)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}>=19'b0001111010010111101) && ({row_reg, col_reg}<19'b0001111010010111111)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0001111010010111111)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0001111010011000000) && ({row_reg, col_reg}<19'b0001111010011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111010011110110) && ({row_reg, col_reg}<19'b0001111010011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111010011111001) && ({row_reg, col_reg}<19'b0001111010100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111010100100001) && ({row_reg, col_reg}<19'b0001111010100100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001111010100100110) && ({row_reg, col_reg}<19'b0001111010100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111010100101001)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==19'b0001111010100101010)) color_data = 12'b110011011000;
		if(({row_reg, col_reg}==19'b0001111010100101011)) color_data = 12'b110111101000;
		if(({row_reg, col_reg}==19'b0001111010100101100)) color_data = 12'b110011010101;
		if(({row_reg, col_reg}==19'b0001111010100101101)) color_data = 12'b110011100101;
		if(({row_reg, col_reg}==19'b0001111010100101110)) color_data = 12'b111011110110;
		if(({row_reg, col_reg}==19'b0001111010100101111)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==19'b0001111010100110000)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0001111010100110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0001111010100110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111010100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001111010100110100) && ({row_reg, col_reg}<19'b0001111010110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111010110000000) && ({row_reg, col_reg}<19'b0001111010110000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001111010110000011) && ({row_reg, col_reg}<19'b0001111010110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111010110000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0001111010110000110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==19'b0001111010110000111)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==19'b0001111010110001000)) color_data = 12'b011000110001;
		if(({row_reg, col_reg}==19'b0001111010110001001)) color_data = 12'b011100110010;
		if(({row_reg, col_reg}==19'b0001111010110001010)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}>=19'b0001111010110001011) && ({row_reg, col_reg}<19'b0001111010110001101)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}==19'b0001111010110001101)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==19'b0001111010110001110)) color_data = 12'b100000100001;
		if(({row_reg, col_reg}==19'b0001111010110001111)) color_data = 12'b011000010001;
		if(({row_reg, col_reg}==19'b0001111010110010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==19'b0001111010110010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111010110010010) && ({row_reg, col_reg}<19'b0001111010110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111010110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111010110011000) && ({row_reg, col_reg}<19'b0001111011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111011001010001) && ({row_reg, col_reg}<19'b0001111011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001111011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001111011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001111100000000000) && ({row_reg, col_reg}<19'b0001111100010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111100010101111)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0001111100010110000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0001111100010110001) && ({row_reg, col_reg}<19'b0001111100010110100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0001111100010110100)) color_data = 12'b001000100110;
		if(({row_reg, col_reg}==19'b0001111100010110101)) color_data = 12'b011001101001;
		if(({row_reg, col_reg}==19'b0001111100010110110)) color_data = 12'b011001011001;
		if(({row_reg, col_reg}==19'b0001111100010110111)) color_data = 12'b010000110110;
		if(({row_reg, col_reg}==19'b0001111100010111000)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}>=19'b0001111100010111001) && ({row_reg, col_reg}<19'b0001111100010111011)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}>=19'b0001111100010111011) && ({row_reg, col_reg}<19'b0001111100010111110)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0001111100010111110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0001111100010111111)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0001111100011000000) && ({row_reg, col_reg}<19'b0001111100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111100011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111100011110001) && ({row_reg, col_reg}<19'b0001111100011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111100011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001111100011110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001111100011110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0001111100011111000) && ({row_reg, col_reg}<19'b0001111100011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111100011111010) && ({row_reg, col_reg}<19'b0001111100100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111100100100001) && ({row_reg, col_reg}<19'b0001111100100100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001111100100100110) && ({row_reg, col_reg}<19'b0001111100100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111100100101001)) color_data = 12'b001100110000;
		if(({row_reg, col_reg}==19'b0001111100100101010)) color_data = 12'b010101010001;
		if(({row_reg, col_reg}==19'b0001111100100101011)) color_data = 12'b011001110001;
		if(({row_reg, col_reg}==19'b0001111100100101100)) color_data = 12'b101010110011;
		if(({row_reg, col_reg}==19'b0001111100100101101)) color_data = 12'b111011110110;
		if(({row_reg, col_reg}==19'b0001111100100101110)) color_data = 12'b111111110110;
		if(({row_reg, col_reg}==19'b0001111100100101111)) color_data = 12'b110111110110;
		if(({row_reg, col_reg}==19'b0001111100100110000)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0001111100100110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001111100100110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0001111100100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001111100100110100) && ({row_reg, col_reg}<19'b0001111100100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111100100110110) && ({row_reg, col_reg}<19'b0001111100110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111100110000000) && ({row_reg, col_reg}<19'b0001111100110000010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001111100110000010) && ({row_reg, col_reg}<19'b0001111100110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111100110000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==19'b0001111100110000110)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==19'b0001111100110000111)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==19'b0001111100110001000)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}>=19'b0001111100110001001) && ({row_reg, col_reg}<19'b0001111100110001011)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}==19'b0001111100110001011)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}==19'b0001111100110001100)) color_data = 12'b100100110011;
		if(({row_reg, col_reg}==19'b0001111100110001101)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==19'b0001111100110001110)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==19'b0001111100110001111)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}==19'b0001111100110010000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==19'b0001111100110010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0001111100110010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111100110010011) && ({row_reg, col_reg}<19'b0001111100110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111100110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111100110011000) && ({row_reg, col_reg}<19'b0001111101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111101001010001) && ({row_reg, col_reg}<19'b0001111101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001111101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001111101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0001111110000000000) && ({row_reg, col_reg}<19'b0001111110010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111110010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111110010110000) && ({row_reg, col_reg}<19'b0001111110010110100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0001111110010110100)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==19'b0001111110010110101)) color_data = 12'b011001011000;
		if(({row_reg, col_reg}==19'b0001111110010110110)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==19'b0001111110010110111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==19'b0001111110010111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001111110010111001)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0001111110010111010) && ({row_reg, col_reg}<19'b0001111110010111101)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0001111110010111101) && ({row_reg, col_reg}<19'b0001111110010111111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0001111110010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001111110011000000) && ({row_reg, col_reg}<19'b0001111110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111110011110000)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0001111110011110001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0001111110011110010) && ({row_reg, col_reg}<19'b0001111110011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111110011110101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==19'b0001111110011110110)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==19'b0001111110011110111)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}>=19'b0001111110011111000) && ({row_reg, col_reg}<19'b0001111110011111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0001111110011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0001111110011111011) && ({row_reg, col_reg}<19'b0001111110100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111110100100010) && ({row_reg, col_reg}<19'b0001111110100100101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0001111110100100101) && ({row_reg, col_reg}<19'b0001111110100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111110100101000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0001111110100101001) && ({row_reg, col_reg}<19'b0001111110100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111110100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0001111110100101100)) color_data = 12'b100010010011;
		if(({row_reg, col_reg}>=19'b0001111110100101101) && ({row_reg, col_reg}<19'b0001111110100101111)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==19'b0001111110100101111)) color_data = 12'b110011010110;
		if(({row_reg, col_reg}==19'b0001111110100110000)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==19'b0001111110100110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0001111110100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001111110100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111110100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0001111110100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0001111110100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111110100110111) && ({row_reg, col_reg}<19'b0001111110101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111110101101010) && ({row_reg, col_reg}<19'b0001111110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111110101101110) && ({row_reg, col_reg}<19'b0001111110101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001111110101110000) && ({row_reg, col_reg}<19'b0001111110110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111110110000000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0001111110110000001) && ({row_reg, col_reg}<19'b0001111110110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111110110000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==19'b0001111110110000110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==19'b0001111110110000111)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==19'b0001111110110001000)) color_data = 12'b101001100110;
		if(({row_reg, col_reg}==19'b0001111110110001001)) color_data = 12'b101001100101;
		if(({row_reg, col_reg}==19'b0001111110110001010)) color_data = 12'b101001010101;
		if(({row_reg, col_reg}==19'b0001111110110001011)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}>=19'b0001111110110001100) && ({row_reg, col_reg}<19'b0001111110110001110)) color_data = 12'b100100110011;
		if(({row_reg, col_reg}==19'b0001111110110001110)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}==19'b0001111110110001111)) color_data = 12'b101001010101;
		if(({row_reg, col_reg}==19'b0001111110110010000)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==19'b0001111110110010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0001111110110010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0001111110110010011) && ({row_reg, col_reg}<19'b0001111110110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0001111110110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0001111110110011000) && ({row_reg, col_reg}<19'b0001111111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0001111111001010001) && ({row_reg, col_reg}<19'b0001111111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0001111111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0001111111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010000000000000000) && ({row_reg, col_reg}<19'b0010000000011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010000000011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000000011000010) && ({row_reg, col_reg}<19'b0010000000011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010000000011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010000000011001000) && ({row_reg, col_reg}<19'b0010000000011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000000011001010) && ({row_reg, col_reg}<19'b0010000000011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000000011011100) && ({row_reg, col_reg}<19'b0010000000011011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010000000011011110) && ({row_reg, col_reg}<19'b0010000000011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000011110001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010000000011110010)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0010000000011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010000000011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010000000011110110)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==19'b0010000000011110111)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==19'b0010000000011111000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==19'b0010000000011111001)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==19'b0010000000011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010000000011111011) && ({row_reg, col_reg}<19'b0010000000100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000100101001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0010000000100101010) && ({row_reg, col_reg}<19'b0010000000100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000100101100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==19'b0010000000100101101)) color_data = 12'b111011101100;
		if(({row_reg, col_reg}==19'b0010000000100101110)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0010000000100101111)) color_data = 12'b110111101011;
		if(({row_reg, col_reg}>=19'b0010000000100110000) && ({row_reg, col_reg}<19'b0010000000110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000000110000110) && ({row_reg, col_reg}<19'b0010000000110001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010000000110001000)) color_data = 12'b011000100011;
		if(({row_reg, col_reg}==19'b0010000000110001001)) color_data = 12'b100001000100;
		if(({row_reg, col_reg}==19'b0010000000110001010)) color_data = 12'b101001010110;
		if(({row_reg, col_reg}==19'b0010000000110001011)) color_data = 12'b101101100111;
		if(({row_reg, col_reg}==19'b0010000000110001100)) color_data = 12'b110001010111;
		if(({row_reg, col_reg}>=19'b0010000000110001101) && ({row_reg, col_reg}<19'b0010000000110001111)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==19'b0010000000110001111)) color_data = 12'b101001010110;
		if(({row_reg, col_reg}==19'b0010000000110010000)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==19'b0010000000110010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010000000110010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010000000110010011) && ({row_reg, col_reg}<19'b0010000000110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000000110011000) && ({row_reg, col_reg}<19'b0010000000110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010000000110111011)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==19'b0010000000110111100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0010000000110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000110111110)) color_data = 12'b011001110011;
		if(({row_reg, col_reg}==19'b0010000000110111111)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==19'b0010000000111000000)) color_data = 12'b100110100110;
		if(({row_reg, col_reg}==19'b0010000000111000001)) color_data = 12'b001101000000;
		if(({row_reg, col_reg}>=19'b0010000000111000010) && ({row_reg, col_reg}<19'b0010000000111000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000000111000111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010000000111001000) && ({row_reg, col_reg}<19'b0010000001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000001001010001) && ({row_reg, col_reg}<19'b0010000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010000001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010000001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010000010000000000) && ({row_reg, col_reg}<19'b0010000010011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000010011000001) && ({row_reg, col_reg}<19'b0010000010011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000010011000100) && ({row_reg, col_reg}<19'b0010000010011001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000010011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000010011001011) && ({row_reg, col_reg}<19'b0010000010011001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010000010011001110) && ({row_reg, col_reg}<19'b0010000010011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000010011010000) && ({row_reg, col_reg}<19'b0010000010011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000010011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010000010011011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010000010011011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010000010011011100) && ({row_reg, col_reg}<19'b0010000010011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000010011011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010000010011100000) && ({row_reg, col_reg}<19'b0010000010011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000010011110001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010000010011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000010011110011) && ({row_reg, col_reg}<19'b0010000010011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000010011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010000010011110110)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==19'b0010000010011110111)) color_data = 12'b100001100011;
		if(({row_reg, col_reg}==19'b0010000010011111000)) color_data = 12'b011001000001;
		if(({row_reg, col_reg}==19'b0010000010011111001)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==19'b0010000010011111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010000010011111011) && ({row_reg, col_reg}<19'b0010000010100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000010100101001) && ({row_reg, col_reg}<19'b0010000010100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010000010100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000010100101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010000010100101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010000010100101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000010100101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0010000010100110000) && ({row_reg, col_reg}<19'b0010000010110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000010110000110) && ({row_reg, col_reg}<19'b0010000010110001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010000010110001000)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0010000010110001001)) color_data = 12'b010100000010;
		if(({row_reg, col_reg}==19'b0010000010110001010)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}==19'b0010000010110001011)) color_data = 12'b100100110101;
		if(({row_reg, col_reg}==19'b0010000010110001100)) color_data = 12'b101000110110;
		if(({row_reg, col_reg}==19'b0010000010110001101)) color_data = 12'b101000110101;
		if(({row_reg, col_reg}==19'b0010000010110001110)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==19'b0010000010110001111)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==19'b0010000010110010000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==19'b0010000010110010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010000010110010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000010110010011) && ({row_reg, col_reg}<19'b0010000010110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000010110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000010110011000) && ({row_reg, col_reg}<19'b0010000010110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000010110110110) && ({row_reg, col_reg}<19'b0010000010110111001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010000010110111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000010110111010) && ({row_reg, col_reg}<19'b0010000010110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010000010110111100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0010000010110111101)) color_data = 12'b001000110000;
		if(({row_reg, col_reg}==19'b0010000010110111110)) color_data = 12'b100110100101;
		if(({row_reg, col_reg}==19'b0010000010110111111)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010000010111000000)) color_data = 12'b101010110110;
		if(({row_reg, col_reg}==19'b0010000010111000001)) color_data = 12'b010001000000;
		if(({row_reg, col_reg}>=19'b0010000010111000010) && ({row_reg, col_reg}<19'b0010000010111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000010111000100)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0010000010111000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000010111000110) && ({row_reg, col_reg}<19'b0010000010111001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000010111001000) && ({row_reg, col_reg}<19'b0010000010111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010000010111001010) && ({row_reg, col_reg}<19'b0010000011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000011001010001) && ({row_reg, col_reg}<19'b0010000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010000011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010000011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010000100000000000) && ({row_reg, col_reg}<19'b0010000100011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000100011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000100011000011) && ({row_reg, col_reg}<19'b0010000100011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000100011000111) && ({row_reg, col_reg}<19'b0010000100011001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010000100011001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010000100011001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000100011001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0010000100011001100) && ({row_reg, col_reg}<19'b0010000100011010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000100011010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010000100011010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000100011010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000100011010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010000100011010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010000100011010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010000100011010111) && ({row_reg, col_reg}<19'b0010000100011011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010000100011011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000100011011100) && ({row_reg, col_reg}<19'b0010000100011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000100011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000100011100000) && ({row_reg, col_reg}<19'b0010000100011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000100011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010000100011110101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010000100011110110)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==19'b0010000100011110111)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==19'b0010000100011111000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==19'b0010000100011111001)) color_data = 12'b010100100000;
		if(({row_reg, col_reg}==19'b0010000100011111010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010000100011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010000100011111100) && ({row_reg, col_reg}<19'b0010000100100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000100100101001) && ({row_reg, col_reg}<19'b0010000100100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010000100100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000100100101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010000100100101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010000100100101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000100100101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010000100100110000) && ({row_reg, col_reg}<19'b0010000100110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000100110000110) && ({row_reg, col_reg}<19'b0010000100110001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010000100110001000) && ({row_reg, col_reg}<19'b0010000100110001010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010000100110001010)) color_data = 12'b010000000001;
		if(({row_reg, col_reg}==19'b0010000100110001011)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}>=19'b0010000100110001100) && ({row_reg, col_reg}<19'b0010000100110001110)) color_data = 12'b100100110101;
		if(({row_reg, col_reg}==19'b0010000100110001110)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==19'b0010000100110001111)) color_data = 12'b010000000001;
		if(({row_reg, col_reg}==19'b0010000100110010000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0010000100110010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000100110010010) && ({row_reg, col_reg}<19'b0010000100110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000100110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000100110011000) && ({row_reg, col_reg}<19'b0010000100110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000100110110110) && ({row_reg, col_reg}<19'b0010000100110111001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010000100110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000100110111010) && ({row_reg, col_reg}<19'b0010000100110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000100110111100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0010000100110111101)) color_data = 12'b011001110011;
		if(({row_reg, col_reg}==19'b0010000100110111110)) color_data = 12'b110111011001;
		if(({row_reg, col_reg}==19'b0010000100110111111)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010000100111000000)) color_data = 12'b110011000111;
		if(({row_reg, col_reg}==19'b0010000100111000001)) color_data = 12'b010101100001;
		if(({row_reg, col_reg}>=19'b0010000100111000010) && ({row_reg, col_reg}<19'b0010000100111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000100111000100) && ({row_reg, col_reg}<19'b0010000100111000110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=19'b0010000100111000110) && ({row_reg, col_reg}<19'b0010000100111001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000100111001000) && ({row_reg, col_reg}<19'b0010000100111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010000100111001010) && ({row_reg, col_reg}<19'b0010000101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000101001010001) && ({row_reg, col_reg}<19'b0010000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010000101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010000101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010000110000000000) && ({row_reg, col_reg}<19'b0010000110011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000110011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000110011000001) && ({row_reg, col_reg}<19'b0010000110011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000110011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010000110011000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010000110011000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000110011000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0010000110011001000) && ({row_reg, col_reg}<19'b0010000110011001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000110011001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010000110011001011) && ({row_reg, col_reg}<19'b0010000110011010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000110011010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010000110011010101) && ({row_reg, col_reg}<19'b0010000110011011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010000110011011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000110011011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010000110011011010) && ({row_reg, col_reg}<19'b0010000110011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000110011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010000110011011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010000110011011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000110011011111) && ({row_reg, col_reg}<19'b0010000110011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000110011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010000110011110101)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010000110011110110)) color_data = 12'b011000110001;
		if(({row_reg, col_reg}==19'b0010000110011110111)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==19'b0010000110011111000)) color_data = 12'b100001000010;
		if(({row_reg, col_reg}==19'b0010000110011111001)) color_data = 12'b010100100000;
		if(({row_reg, col_reg}==19'b0010000110011111010)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010000110011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010000110011111100) && ({row_reg, col_reg}<19'b0010000110100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000110100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000110100101101) && ({row_reg, col_reg}<19'b0010000110100101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010000110100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000110100110000) && ({row_reg, col_reg}<19'b0010000110110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000110110000110) && ({row_reg, col_reg}<19'b0010000110110001000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010000110110001000) && ({row_reg, col_reg}<19'b0010000110110001010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010000110110001010)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010000110110001011)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==19'b0010000110110001100)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==19'b0010000110110001101)) color_data = 12'b101001010111;
		if(({row_reg, col_reg}==19'b0010000110110001110)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==19'b0010000110110001111)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010000110110010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010000110110010001) && ({row_reg, col_reg}<19'b0010000110110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000110110110110) && ({row_reg, col_reg}<19'b0010000110110111001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010000110110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010000110110111010) && ({row_reg, col_reg}<19'b0010000110110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010000110110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010000110110111101)) color_data = 12'b101010110111;
		if(({row_reg, col_reg}==19'b0010000110110111110)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}>=19'b0010000110110111111) && ({row_reg, col_reg}<19'b0010000110111000001)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==19'b0010000110111000001)) color_data = 12'b011001110010;
		if(({row_reg, col_reg}>=19'b0010000110111000010) && ({row_reg, col_reg}<19'b0010000110111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000110111000100) && ({row_reg, col_reg}<19'b0010000110111000110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0010000110111000110) && ({row_reg, col_reg}<19'b0010000110111001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000110111001000) && ({row_reg, col_reg}<19'b0010000110111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010000110111001010) && ({row_reg, col_reg}<19'b0010000111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010000111001010001) && ({row_reg, col_reg}<19'b0010000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010000111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010000111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010001000000000000) && ({row_reg, col_reg}<19'b0010001000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001000011000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010001000011000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0010001000011000101) && ({row_reg, col_reg}<19'b0010001000011001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001000011001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001000011001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001000011001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000011001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010001000011001110) && ({row_reg, col_reg}<19'b0010001000011010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010001000011010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010001000011010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000011010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001000011010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001000011010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010001000011010110) && ({row_reg, col_reg}<19'b0010001000011011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001000011011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010001000011011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010001000011011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010001000011011100) && ({row_reg, col_reg}<19'b0010001000011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010001000011011111) && ({row_reg, col_reg}<19'b0010001000011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001000011110010) && ({row_reg, col_reg}<19'b0010001000011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010001000011110100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010001000011110101)) color_data = 12'b010100010000;
		if(({row_reg, col_reg}==19'b0010001000011110110)) color_data = 12'b100001000010;
		if(({row_reg, col_reg}==19'b0010001000011110111)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}==19'b0010001000011111000)) color_data = 12'b100101000010;
		if(({row_reg, col_reg}==19'b0010001000011111001)) color_data = 12'b011100110001;
		if(({row_reg, col_reg}==19'b0010001000011111010)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==19'b0010001000011111011)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010001000011111100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010001000011111101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0010001000011111110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0010001000011111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010001000100000000) && ({row_reg, col_reg}<19'b0010001000100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001000100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010001000100101110) && ({row_reg, col_reg}<19'b0010001000110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001000110000111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010001000110001000) && ({row_reg, col_reg}<19'b0010001000110001010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010001000110001010)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010001000110001011)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==19'b0010001000110001100)) color_data = 12'b100101000110;
		if(({row_reg, col_reg}==19'b0010001000110001101)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==19'b0010001000110001110)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==19'b0010001000110001111)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}>=19'b0010001000110010000) && ({row_reg, col_reg}<19'b0010001000110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001000110110110) && ({row_reg, col_reg}<19'b0010001000110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010001000110111000) && ({row_reg, col_reg}<19'b0010001000110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001000110111100)) color_data = 12'b001101000001;
		if(({row_reg, col_reg}==19'b0010001000110111101)) color_data = 12'b110011011001;
		if(({row_reg, col_reg}==19'b0010001000110111110)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==19'b0010001000110111111)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0010001000111000000)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010001000111000001)) color_data = 12'b100010010101;
		if(({row_reg, col_reg}==19'b0010001000111000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=19'b0010001000111000011) && ({row_reg, col_reg}<19'b0010001000111001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001000111001000) && ({row_reg, col_reg}<19'b0010001000111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010001000111001010) && ({row_reg, col_reg}<19'b0010001001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001001001010001) && ({row_reg, col_reg}<19'b0010001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010001001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010001001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010001010000000000) && ({row_reg, col_reg}<19'b0010001010010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001010010111110) && ({row_reg, col_reg}<19'b0010001010011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010001010011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001010011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010001010011000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010001010011000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0010001010011000100) && ({row_reg, col_reg}<19'b0010001010011000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001010011000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010001010011000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001010011001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010011001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010001010011001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010001010011001011) && ({row_reg, col_reg}<19'b0010001010011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001010011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010001010011010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010001010011010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010001010011010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010001010011010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010011010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001010011011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010001010011011001) && ({row_reg, col_reg}<19'b0010001010011011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001010011011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001010011011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010001010011011101) && ({row_reg, col_reg}<19'b0010001010011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001010011011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010001010011100000) && ({row_reg, col_reg}<19'b0010001010011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001010011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010001010011110010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010001010011110011)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010001010011110100)) color_data = 12'b010100010001;
		if(({row_reg, col_reg}==19'b0010001010011110101)) color_data = 12'b011100100010;
		if(({row_reg, col_reg}==19'b0010001010011110110)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}==19'b0010001010011110111)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}==19'b0010001010011111000)) color_data = 12'b100101000010;
		if(({row_reg, col_reg}==19'b0010001010011111001)) color_data = 12'b100000110010;
		if(({row_reg, col_reg}==19'b0010001010011111010)) color_data = 12'b011000100001;
		if(({row_reg, col_reg}==19'b0010001010011111011)) color_data = 12'b010100100001;
		if(({row_reg, col_reg}==19'b0010001010011111100)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==19'b0010001010011111101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==19'b0010001010011111110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0010001010011111111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0010001010100000000) && ({row_reg, col_reg}<19'b0010001010110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001010110000111) && ({row_reg, col_reg}<19'b0010001010110001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010001010110001010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010001010110001011)) color_data = 12'b010000000001;
		if(({row_reg, col_reg}==19'b0010001010110001100)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==19'b0010001010110001101)) color_data = 12'b011000100011;
		if(({row_reg, col_reg}==19'b0010001010110001110)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==19'b0010001010110001111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0010001010110010000) && ({row_reg, col_reg}<19'b0010001010110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001010110110110) && ({row_reg, col_reg}<19'b0010001010110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010001010110111000) && ({row_reg, col_reg}<19'b0010001010110111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001010110111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0010001010110111100)) color_data = 12'b100010000101;
		if(({row_reg, col_reg}==19'b0010001010110111101)) color_data = 12'b110111101010;
		if(({row_reg, col_reg}==19'b0010001010110111110)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010001010110111111)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0010001010111000000)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010001010111000001)) color_data = 12'b101111000111;
		if(({row_reg, col_reg}==19'b0010001010111000010)) color_data = 12'b011001110011;
		if(({row_reg, col_reg}==19'b0010001010111000011)) color_data = 12'b010001000001;
		if(({row_reg, col_reg}==19'b0010001010111000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=19'b0010001010111000101) && ({row_reg, col_reg}<19'b0010001010111000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001010111000111) && ({row_reg, col_reg}<19'b0010001010111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010001010111001010) && ({row_reg, col_reg}<19'b0010001011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001011001010001) && ({row_reg, col_reg}<19'b0010001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010001011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010001011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010001100000000000) && ({row_reg, col_reg}<19'b0010001100010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001100010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010001100010111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010001100011000000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010001100011000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001100011000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001100011000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010001100011000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010001100011000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001100011000110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010001100011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010001100011001000) && ({row_reg, col_reg}<19'b0010001100011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001100011001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010001100011001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010001100011010000) && ({row_reg, col_reg}<19'b0010001100011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010001100011010100) && ({row_reg, col_reg}<19'b0010001100011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001100011011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010001100011011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0010001100011011010) && ({row_reg, col_reg}<19'b0010001100011011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001100011011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001100011011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010001100011011110) && ({row_reg, col_reg}<19'b0010001100011100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010001100011100000) && ({row_reg, col_reg}<19'b0010001100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001100011110000) && ({row_reg, col_reg}<19'b0010001100011110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010001100011110010)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0010001100011110011)) color_data = 12'b010100010010;
		if(({row_reg, col_reg}==19'b0010001100011110100)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}==19'b0010001100011110101)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}>=19'b0010001100011110110) && ({row_reg, col_reg}<19'b0010001100011111000)) color_data = 12'b101001000011;
		if(({row_reg, col_reg}==19'b0010001100011111000)) color_data = 12'b100101000010;
		if(({row_reg, col_reg}==19'b0010001100011111001)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==19'b0010001100011111010)) color_data = 12'b100000110011;
		if(({row_reg, col_reg}==19'b0010001100011111011)) color_data = 12'b100001000100;
		if(({row_reg, col_reg}==19'b0010001100011111100)) color_data = 12'b100001000101;
		if(({row_reg, col_reg}==19'b0010001100011111101)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==19'b0010001100011111110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0010001100011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010001100100000000) && ({row_reg, col_reg}<19'b0010001100110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001100110000111) && ({row_reg, col_reg}<19'b0010001100110001001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010001100110001001) && ({row_reg, col_reg}<19'b0010001100110001011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010001100110001011)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}>=19'b0010001100110001100) && ({row_reg, col_reg}<19'b0010001100110001110)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0010001100110001110)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010001100110001111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010001100110010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010001100110010001) && ({row_reg, col_reg}<19'b0010001100110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001100110110110) && ({row_reg, col_reg}<19'b0010001100110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010001100110111000) && ({row_reg, col_reg}<19'b0010001100110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001100110111010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==19'b0010001100110111011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==19'b0010001100110111100)) color_data = 12'b110111011010;
		if(({row_reg, col_reg}==19'b0010001100110111101)) color_data = 12'b111011111011;
		if(({row_reg, col_reg}>=19'b0010001100110111110) && ({row_reg, col_reg}<19'b0010001100111000000)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==19'b0010001100111000000)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==19'b0010001100111000001)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0010001100111000010)) color_data = 12'b110011011001;
		if(({row_reg, col_reg}==19'b0010001100111000011)) color_data = 12'b101010111000;
		if(({row_reg, col_reg}==19'b0010001100111000100)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==19'b0010001100111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010001100111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001100111000111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0010001100111001000) && ({row_reg, col_reg}<19'b0010001100111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010001100111001010) && ({row_reg, col_reg}<19'b0010001101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001101001010001) && ({row_reg, col_reg}<19'b0010001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010001101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010001101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010001110000000000) && ({row_reg, col_reg}<19'b0010001110010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001110010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010001110010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010001110010111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010001110011000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010001110011000001) && ({row_reg, col_reg}<19'b0010001110011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001110011000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001110011000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010001110011000101) && ({row_reg, col_reg}<19'b0010001110011011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001110011011010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010001110011011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0010001110011011100) && ({row_reg, col_reg}<19'b0010001110011011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001110011011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010001110011011111) && ({row_reg, col_reg}<19'b0010001110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001110011110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010001110011110001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010001110011110010)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0010001110011110011)) color_data = 12'b011000100011;
		if(({row_reg, col_reg}==19'b0010001110011110100)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==19'b0010001110011110101)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}==19'b0010001110011110110)) color_data = 12'b101101010100;
		if(({row_reg, col_reg}==19'b0010001110011110111)) color_data = 12'b101001000011;
		if(({row_reg, col_reg}==19'b0010001110011111000)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==19'b0010001110011111001)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}==19'b0010001110011111010)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==19'b0010001110011111011)) color_data = 12'b101001010101;
		if(({row_reg, col_reg}==19'b0010001110011111100)) color_data = 12'b100101010110;
		if(({row_reg, col_reg}==19'b0010001110011111101)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==19'b0010001110011111110)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==19'b0010001110011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010001110100000000) && ({row_reg, col_reg}<19'b0010001110110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001110110001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0010001110110001001) && ({row_reg, col_reg}<19'b0010001110110001011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0010001110110001011)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}>=19'b0010001110110001100) && ({row_reg, col_reg}<19'b0010001110110001110)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010001110110001110)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010001110110001111)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0010001110110010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010001110110010001) && ({row_reg, col_reg}<19'b0010001110110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010001110110010101) && ({row_reg, col_reg}<19'b0010001110110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001110110110110) && ({row_reg, col_reg}<19'b0010001110110111001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010001110110111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010001110110111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010001110110111011)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}==19'b0010001110110111100)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0010001110110111101)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010001110110111110)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0010001110110111111)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010001110111000000)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0010001110111000001)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010001110111000010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==19'b0010001110111000011)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0010001110111000100)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==19'b0010001110111000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==19'b0010001110111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001110111000111) && ({row_reg, col_reg}<19'b0010001110111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010001110111001010) && ({row_reg, col_reg}<19'b0010001111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010001111001010001) && ({row_reg, col_reg}<19'b0010001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010001111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010001111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010010000000000000) && ({row_reg, col_reg}<19'b0010010000010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010000010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010010000010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010010000010110011) && ({row_reg, col_reg}<19'b0010010000010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010000010111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010010000010111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0010010000010111111) && ({row_reg, col_reg}<19'b0010010000011000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010000011000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010000011000010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010010000011000011) && ({row_reg, col_reg}<19'b0010010000011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010000011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010000011000110) && ({row_reg, col_reg}<19'b0010010000011010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010000011010001) && ({row_reg, col_reg}<19'b0010010000011010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010010000011010011) && ({row_reg, col_reg}<19'b0010010000011010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010000011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010000011010110) && ({row_reg, col_reg}<19'b0010010000011011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010010000011011000) && ({row_reg, col_reg}<19'b0010010000011011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010000011011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010010000011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010010000011011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010000011011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010000011011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010010000011011111) && ({row_reg, col_reg}<19'b0010010000011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010000011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010010000011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010010000011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010000011100100) && ({row_reg, col_reg}<19'b0010010000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010000011110000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0010010000011110001)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0010010000011110010)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==19'b0010010000011110011)) color_data = 12'b011000100010;
		if(({row_reg, col_reg}==19'b0010010000011110100)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}==19'b0010010000011110101)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}==19'b0010010000011110110)) color_data = 12'b101001000011;
		if(({row_reg, col_reg}>=19'b0010010000011110111) && ({row_reg, col_reg}<19'b0010010000011111001)) color_data = 12'b101101010100;
		if(({row_reg, col_reg}==19'b0010010000011111001)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}==19'b0010010000011111010)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==19'b0010010000011111011)) color_data = 12'b100001000100;
		if(({row_reg, col_reg}==19'b0010010000011111100)) color_data = 12'b011000100011;
		if(({row_reg, col_reg}==19'b0010010000011111101)) color_data = 12'b010100010010;
		if(({row_reg, col_reg}==19'b0010010000011111110)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0010010000011111111)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0010010000100000000) && ({row_reg, col_reg}<19'b0010010000110001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010000110001001) && ({row_reg, col_reg}<19'b0010010000110010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010010000110010000) && ({row_reg, col_reg}<19'b0010010000110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010000110110110) && ({row_reg, col_reg}<19'b0010010000110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010010000110111000) && ({row_reg, col_reg}<19'b0010010000110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010000110111010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==19'b0010010000110111011)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==19'b0010010000110111100)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0010010000110111101)) color_data = 12'b101110110111;
		if(({row_reg, col_reg}==19'b0010010000110111110)) color_data = 12'b101111000111;
		if(({row_reg, col_reg}==19'b0010010000110111111)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010010000111000000)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}>=19'b0010010000111000001) && ({row_reg, col_reg}<19'b0010010000111000011)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==19'b0010010000111000011)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==19'b0010010000111000100)) color_data = 12'b010101100100;
		if(({row_reg, col_reg}==19'b0010010000111000101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==19'b0010010000111000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010010000111000111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0010010000111001000) && ({row_reg, col_reg}<19'b0010010000111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010010000111001010) && ({row_reg, col_reg}<19'b0010010001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010001001010001) && ({row_reg, col_reg}<19'b0010010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010010001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010010001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010010010000000000) && ({row_reg, col_reg}<19'b0010010010010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010010010110001) && ({row_reg, col_reg}<19'b0010010010010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010010010110011) && ({row_reg, col_reg}<19'b0010010010010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010010010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010010010010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010010010010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010010010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010010010111001) && ({row_reg, col_reg}<19'b0010010010010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010010010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010010010010111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010010010010111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010010010111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010010010010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010010011000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010010010011000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010010010011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010010011000011) && ({row_reg, col_reg}<19'b0010010010011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010010011000101) && ({row_reg, col_reg}<19'b0010010010011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010010011001000) && ({row_reg, col_reg}<19'b0010010010011001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010010011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010010010011001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010010010011001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010010010011001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010010010011001110) && ({row_reg, col_reg}<19'b0010010010011010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010010011010001) && ({row_reg, col_reg}<19'b0010010010011010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010010011010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010010010011010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010010010011010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010010010011010110) && ({row_reg, col_reg}<19'b0010010010011011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010010011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010010010011011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010010010011011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010010011011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010010011011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010010010011011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010010010011100000) && ({row_reg, col_reg}<19'b0010010010011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010010011100010) && ({row_reg, col_reg}<19'b0010010010011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010010011100100) && ({row_reg, col_reg}<19'b0010010010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010010011110000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0010010010011110001)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0010010010011110010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010010010011110011)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010010010011110100)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==19'b0010010010011110101)) color_data = 12'b010100000000;
		if(({row_reg, col_reg}==19'b0010010010011110110)) color_data = 12'b011000010000;
		if(({row_reg, col_reg}==19'b0010010010011110111)) color_data = 12'b011100010000;
		if(({row_reg, col_reg}==19'b0010010010011111000)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==19'b0010010010011111001)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}==19'b0010010010011111010)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==19'b0010010010011111011)) color_data = 12'b100000110011;
		if(({row_reg, col_reg}==19'b0010010010011111100)) color_data = 12'b010100010010;
		if(({row_reg, col_reg}==19'b0010010010011111101)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}>=19'b0010010010011111110) && ({row_reg, col_reg}<19'b0010010010100000000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0010010010100000000) && ({row_reg, col_reg}<19'b0010010010110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010010110001100) && ({row_reg, col_reg}<19'b0010010010110001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010010010110001111) && ({row_reg, col_reg}<19'b0010010010110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010010110110110) && ({row_reg, col_reg}<19'b0010010010110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010010010110111000) && ({row_reg, col_reg}<19'b0010010010110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010010110111010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}>=19'b0010010010110111011) && ({row_reg, col_reg}<19'b0010010010110111101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==19'b0010010010110111101)) color_data = 12'b010101010010;
		if(({row_reg, col_reg}==19'b0010010010110111110)) color_data = 12'b011101110011;
		if(({row_reg, col_reg}==19'b0010010010110111111)) color_data = 12'b110011011000;
		if(({row_reg, col_reg}==19'b0010010010111000000)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0010010010111000001)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==19'b0010010010111000010)) color_data = 12'b110011011001;
		if(({row_reg, col_reg}==19'b0010010010111000011)) color_data = 12'b011101110100;
		if(({row_reg, col_reg}==19'b0010010010111000100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0010010010111000101) && ({row_reg, col_reg}<19'b0010010010111001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010010111001000) && ({row_reg, col_reg}<19'b0010010010111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010010010111001010) && ({row_reg, col_reg}<19'b0010010011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010011001010001) && ({row_reg, col_reg}<19'b0010010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010010011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010010011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010010100000000000) && ({row_reg, col_reg}<19'b0010010100010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010100010110000) && ({row_reg, col_reg}<19'b0010010100010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010100010110010) && ({row_reg, col_reg}<19'b0010010100010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010100010110101) && ({row_reg, col_reg}<19'b0010010100010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010010100010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010100010111000) && ({row_reg, col_reg}<19'b0010010100010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010100010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010010100010111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010100010111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010010100010111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010100010111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010100010111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010100011000000) && ({row_reg, col_reg}<19'b0010010100011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010100011000011) && ({row_reg, col_reg}<19'b0010010100011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010100011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010010100011001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010010100011001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010010100011001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010100011001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010100011001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010010100011001101) && ({row_reg, col_reg}<19'b0010010100011010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010100011010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010010100011010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010100011010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010010100011010111) && ({row_reg, col_reg}<19'b0010010100011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010100011011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010010100011011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010010100011011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010100011011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010100011011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0010010100011100000) && ({row_reg, col_reg}<19'b0010010100011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010100011100011) && ({row_reg, col_reg}<19'b0010010100011100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010100011100101) && ({row_reg, col_reg}<19'b0010010100011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010100011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010100011101000) && ({row_reg, col_reg}<19'b0010010100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010100011110000) && ({row_reg, col_reg}<19'b0010010100011110010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0010010100011110010) && ({row_reg, col_reg}<19'b0010010100011110101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0010010100011110101) && ({row_reg, col_reg}<19'b0010010100011111000)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010010100011111000)) color_data = 12'b011000010000;
		if(({row_reg, col_reg}==19'b0010010100011111001)) color_data = 12'b100000110010;
		if(({row_reg, col_reg}==19'b0010010100011111010)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==19'b0010010100011111011)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}==19'b0010010100011111100)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}>=19'b0010010100011111101) && ({row_reg, col_reg}<19'b0010010100011111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010010100011111111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=19'b0010010100100000000) && ({row_reg, col_reg}<19'b0010010100110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010100110110110) && ({row_reg, col_reg}<19'b0010010100110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010010100110111000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0010010100110111001) && ({row_reg, col_reg}<19'b0010010100110111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010100110111011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0010010100110111100)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0010010100110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010100110111110)) color_data = 12'b001101000000;
		if(({row_reg, col_reg}==19'b0010010100110111111)) color_data = 12'b100110010100;
		if(({row_reg, col_reg}==19'b0010010100111000000)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==19'b0010010100111000001)) color_data = 12'b110111101010;
		if(({row_reg, col_reg}==19'b0010010100111000010)) color_data = 12'b100110100110;
		if(({row_reg, col_reg}==19'b0010010100111000011)) color_data = 12'b001101000001;
		if(({row_reg, col_reg}>=19'b0010010100111000100) && ({row_reg, col_reg}<19'b0010010100111001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010100111001000) && ({row_reg, col_reg}<19'b0010010100111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010010100111001010) && ({row_reg, col_reg}<19'b0010010101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010101001010001) && ({row_reg, col_reg}<19'b0010010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010010101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010010101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010010110000000000) && ({row_reg, col_reg}<19'b0010010110010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010110010110000) && ({row_reg, col_reg}<19'b0010010110010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010110010110010) && ({row_reg, col_reg}<19'b0010010110010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010110010110101) && ({row_reg, col_reg}<19'b0010010110010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010110010110111) && ({row_reg, col_reg}<19'b0010010110010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010110010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010010110010111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010110010111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010010110010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010110010111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010110010111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010010110010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010110011000000) && ({row_reg, col_reg}<19'b0010010110011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010010110011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010110011000011) && ({row_reg, col_reg}<19'b0010010110011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010110011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010010110011000110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010010110011000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010110011001000) && ({row_reg, col_reg}<19'b0010010110011001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010110011001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010010110011001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010010110011001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010110011001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010110011010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010110011010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010110011010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010110011010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010010110011010100) && ({row_reg, col_reg}<19'b0010010110011010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010110011010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010010110011010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010110011011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010010110011011001) && ({row_reg, col_reg}<19'b0010010110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010110011011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010010110011011110) && ({row_reg, col_reg}<19'b0010010110011100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010010110011100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010010110011100001) && ({row_reg, col_reg}<19'b0010010110011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010110011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010110011100101) && ({row_reg, col_reg}<19'b0010010110011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010110011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010010110011101000) && ({row_reg, col_reg}<19'b0010010110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010110011110000) && ({row_reg, col_reg}<19'b0010010110011110010)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0010010110011110010)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0010010110011110011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0010010110011110100) && ({row_reg, col_reg}<19'b0010010110011111000)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010010110011111000)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==19'b0010010110011111001)) color_data = 12'b011100110001;
		if(({row_reg, col_reg}==19'b0010010110011111010)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==19'b0010010110011111011)) color_data = 12'b011000110011;
		if(({row_reg, col_reg}==19'b0010010110011111100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010010110011111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010010110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010110011111111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0010010110100000000) && ({row_reg, col_reg}<19'b0010010110110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010110110110110) && ({row_reg, col_reg}<19'b0010010110110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010010110110111000)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0010010110110111001) && ({row_reg, col_reg}<19'b0010010110110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010110110111110)) color_data = 12'b001000110000;
		if(({row_reg, col_reg}==19'b0010010110110111111)) color_data = 12'b011110000011;
		if(({row_reg, col_reg}==19'b0010010110111000000)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010010110111000001)) color_data = 12'b110011011001;
		if(({row_reg, col_reg}==19'b0010010110111000010)) color_data = 12'b011101110011;
		if(({row_reg, col_reg}==19'b0010010110111000011)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0010010110111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010010110111000101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==19'b0010010110111000110)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==19'b0010010110111000111)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0010010110111001000) && ({row_reg, col_reg}<19'b0010010110111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010010110111001010) && ({row_reg, col_reg}<19'b0010010111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010010111001010001) && ({row_reg, col_reg}<19'b0010010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010010111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010010111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010011000000000000) && ({row_reg, col_reg}<19'b0010011000010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011000010110001) && ({row_reg, col_reg}<19'b0010011000010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011000010110011) && ({row_reg, col_reg}<19'b0010011000010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011000010110101) && ({row_reg, col_reg}<19'b0010011000010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000010111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010011000010111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0010011000010111010) && ({row_reg, col_reg}<19'b0010011000010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011000010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011000010111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010011000010111110) && ({row_reg, col_reg}<19'b0010011000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000011000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010011000011000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011000011000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011000011000110) && ({row_reg, col_reg}<19'b0010011000011001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011000011001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010011000011001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010011000011001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011000011001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000011001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010011000011001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010011000011001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011000011001111) && ({row_reg, col_reg}<19'b0010011000011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011000011010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011000011010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010011000011010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000011010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011000011010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010011000011010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011000011011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011000011011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011000011011010) && ({row_reg, col_reg}<19'b0010011000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000011011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010011000011011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011000011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011000011100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010011000011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011000011100010) && ({row_reg, col_reg}<19'b0010011000011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011000011100101) && ({row_reg, col_reg}<19'b0010011000011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000011100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011000011101000) && ({row_reg, col_reg}<19'b0010011000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011000011110000) && ({row_reg, col_reg}<19'b0010011000011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011000011110011) && ({row_reg, col_reg}<19'b0010011000011110101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0010011000011110101) && ({row_reg, col_reg}<19'b0010011000011110111)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010011000011110111)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==19'b0010011000011111000)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010011000011111001)) color_data = 12'b011000100001;
		if(({row_reg, col_reg}==19'b0010011000011111010)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==19'b0010011000011111011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==19'b0010011000011111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010011000011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000011111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010011000011111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010011000100000000) && ({row_reg, col_reg}<19'b0010011000110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011000110110110) && ({row_reg, col_reg}<19'b0010011000110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010011000110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011000110111001) && ({row_reg, col_reg}<19'b0010011000110111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000110111011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0010011000110111100) && ({row_reg, col_reg}<19'b0010011000110111110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010011000110111110)) color_data = 12'b001000110000;
		if(({row_reg, col_reg}==19'b0010011000110111111)) color_data = 12'b010101100001;
		if(({row_reg, col_reg}==19'b0010011000111000000)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010011000111000001)) color_data = 12'b101111000111;
		if(({row_reg, col_reg}==19'b0010011000111000010)) color_data = 12'b010101010001;
		if(({row_reg, col_reg}>=19'b0010011000111000011) && ({row_reg, col_reg}<19'b0010011000111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011000111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010011000111000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011000111000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011000111001000) && ({row_reg, col_reg}<19'b0010011000111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010011000111001010) && ({row_reg, col_reg}<19'b0010011001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011001001010001) && ({row_reg, col_reg}<19'b0010011001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010011001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010011001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010011010000000000) && ({row_reg, col_reg}<19'b0010011010010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011010010110011) && ({row_reg, col_reg}<19'b0010011010010110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011010010110101) && ({row_reg, col_reg}<19'b0010011010010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010011010010111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011010010111001) && ({row_reg, col_reg}<19'b0010011010010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011010010111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011010010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011010010111101) && ({row_reg, col_reg}<19'b0010011010010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011010011000000) && ({row_reg, col_reg}<19'b0010011010011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010011000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010011010011000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0010011010011000100) && ({row_reg, col_reg}<19'b0010011010011000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011010011000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010011010011000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011010011001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010011010011001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010011010011001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011010011001011) && ({row_reg, col_reg}<19'b0010011010011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011010011010001) && ({row_reg, col_reg}<19'b0010011010011010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010011010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010011010011010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011010011010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011010011011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010011010011011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010011010011011010) && ({row_reg, col_reg}<19'b0010011010011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011010011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010011011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011010011011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011010011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011010011100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011010011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011010011100010) && ({row_reg, col_reg}<19'b0010011010011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011010011100101) && ({row_reg, col_reg}<19'b0010011010011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010011100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011010011101000) && ({row_reg, col_reg}<19'b0010011010011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010011010011110101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0010011010011110110) && ({row_reg, col_reg}<19'b0010011010011111000)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0010011010011111000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010011010011111001)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==19'b0010011010011111010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==19'b0010011010011111011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==19'b0010011010011111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010011010011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010011111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010011010011111111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0010011010100000000) && ({row_reg, col_reg}<19'b0010011010110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011010110110110) && ({row_reg, col_reg}<19'b0010011010110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010011010110111000) && ({row_reg, col_reg}<19'b0010011010110111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011010110111011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0010011010110111100)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010011010110111101)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0010011010110111110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0010011010110111111)) color_data = 12'b001000110000;
		if(({row_reg, col_reg}==19'b0010011010111000000)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0010011010111000001)) color_data = 12'b110011011000;
		if(({row_reg, col_reg}==19'b0010011010111000010)) color_data = 12'b011001110011;
		if(({row_reg, col_reg}==19'b0010011010111000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0010011010111000100) && ({row_reg, col_reg}<19'b0010011010111001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011010111001000) && ({row_reg, col_reg}<19'b0010011010111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010011010111001010) && ({row_reg, col_reg}<19'b0010011011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011011001010001) && ({row_reg, col_reg}<19'b0010011011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010011011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010011011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010011100000000000) && ({row_reg, col_reg}<19'b0010011100010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011100010110010) && ({row_reg, col_reg}<19'b0010011100010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011100010110100) && ({row_reg, col_reg}<19'b0010011100010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100010110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010011100010110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011100010111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011100010111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010011100010111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011100010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011100010111100) && ({row_reg, col_reg}<19'b0010011100010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010011100011000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010011100011000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011100011000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010011100011000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010011100011000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010011100011000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011100011000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010011100011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011100011001000) && ({row_reg, col_reg}<19'b0010011100011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100011001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011100011010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010011100011010001) && ({row_reg, col_reg}<19'b0010011100011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011100011010100) && ({row_reg, col_reg}<19'b0010011100011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100011010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010011100011010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010011100011011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011100011011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010011100011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011100011011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010011100011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100011011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011100011011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011100011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011100011100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011100011100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011100011100010) && ({row_reg, col_reg}<19'b0010011100011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011100011100101) && ({row_reg, col_reg}<19'b0010011100011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011100011101000) && ({row_reg, col_reg}<19'b0010011100011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011100011110101) && ({row_reg, col_reg}<19'b0010011100011110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010011100011110111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010011100011111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0010011100011111001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0010011100011111010)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==19'b0010011100011111011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=19'b0010011100011111100) && ({row_reg, col_reg}<19'b0010011100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100011111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010011100011111111)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0010011100100000000) && ({row_reg, col_reg}<19'b0010011100110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011100110110110) && ({row_reg, col_reg}<19'b0010011100110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010011100110111000) && ({row_reg, col_reg}<19'b0010011100110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100110111100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0010011100110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010011100110111110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0010011100110111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100111000000)) color_data = 12'b101110110110;
		if(({row_reg, col_reg}==19'b0010011100111000001)) color_data = 12'b101010100110;
		if(({row_reg, col_reg}==19'b0010011100111000010)) color_data = 12'b011001110011;
		if(({row_reg, col_reg}==19'b0010011100111000011)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0010011100111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011100111000101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010011100111000110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0010011100111000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011100111001000) && ({row_reg, col_reg}<19'b0010011100111001010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0010011100111001010) && ({row_reg, col_reg}<19'b0010011101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011101001010001) && ({row_reg, col_reg}<19'b0010011101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010011101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010011101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010011110000000000) && ({row_reg, col_reg}<19'b0010011110010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011110010110001) && ({row_reg, col_reg}<19'b0010011110010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011110010110100) && ({row_reg, col_reg}<19'b0010011110010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110010110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011110010110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011110010111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010011110010111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010011110010111010) && ({row_reg, col_reg}<19'b0010011110010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011110010111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010011110010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011110010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110011000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011110011000001) && ({row_reg, col_reg}<19'b0010011110011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011110011000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011110011000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010011110011000101) && ({row_reg, col_reg}<19'b0010011110011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011110011010010) && ({row_reg, col_reg}<19'b0010011110011010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010011110011010100) && ({row_reg, col_reg}<19'b0010011110011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110011010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010011110011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011110011011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011110011011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010011110011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011110011011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010011110011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110011011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010011110011011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011110011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011110011100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011110011100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010011110011100010) && ({row_reg, col_reg}<19'b0010011110011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011110011100101) && ({row_reg, col_reg}<19'b0010011110011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010011110011101000) && ({row_reg, col_reg}<19'b0010011110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011110011110000) && ({row_reg, col_reg}<19'b0010011110011110011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0010011110011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011110011110100) && ({row_reg, col_reg}<19'b0010011110011111011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0010011110011111011) && ({row_reg, col_reg}<19'b0010011110110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110110111000)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0010011110110111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010011110110111010)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0010011110110111011) && ({row_reg, col_reg}<19'b0010011110110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110110111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0010011110110111110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0010011110110111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010011110111000000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0010011110111000001)) color_data = 12'b001100110000;
		if(({row_reg, col_reg}==19'b0010011110111000010)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}>=19'b0010011110111000011) && ({row_reg, col_reg}<19'b0010011111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010011111001010001) && ({row_reg, col_reg}<19'b0010011111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010011111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010011111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010100000000000000) && ({row_reg, col_reg}<19'b0010100000010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000010110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010100000010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100000010110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100000010111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100000010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100000010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100000010111011) && ({row_reg, col_reg}<19'b0010100000010111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010100000010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010100000010111111) && ({row_reg, col_reg}<19'b0010100000011000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100000011000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100000011000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010100000011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100000011000100) && ({row_reg, col_reg}<19'b0010100000011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000011010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010100000011010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010100000011011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100000011011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0010100000011011010) && ({row_reg, col_reg}<19'b0010100000011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100000011011100) && ({row_reg, col_reg}<19'b0010100000011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000011011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100000011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100000011100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100000011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100000011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100000011100100) && ({row_reg, col_reg}<19'b0010100000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100000100100110) && ({row_reg, col_reg}<19'b0010100000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000100101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010100000100101001) && ({row_reg, col_reg}<19'b0010100000100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100000100101011) && ({row_reg, col_reg}<19'b0010100000100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100000100101101) && ({row_reg, col_reg}<19'b0010100000100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010100000100110000) && ({row_reg, col_reg}<19'b0010100000100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100000100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100000100111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010100000100111100) && ({row_reg, col_reg}<19'b0010100000101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100000101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100000101000001) && ({row_reg, col_reg}<19'b0010100000101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100000101000011) && ({row_reg, col_reg}<19'b0010100000101000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010100000101000101) && ({row_reg, col_reg}<19'b0010100001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100001001010001) && ({row_reg, col_reg}<19'b0010100001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010100001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010100001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010100010000000000) && ({row_reg, col_reg}<19'b0010100010010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100010010110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010100010010110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100010010110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100010010111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010100010010111001) && ({row_reg, col_reg}<19'b0010100010010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010010111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010100010010111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010010111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100010010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100010011000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100010011000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010100010011000011) && ({row_reg, col_reg}<19'b0010100010011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010011010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010100010011010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010100010011011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010100010011011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100010011011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010100010011011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010100010011011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010100010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010011011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100010011011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010100010011100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100010011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100010011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100010011100100) && ({row_reg, col_reg}<19'b0010100010100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010100010100110000) && ({row_reg, col_reg}<19'b0010100010100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100010100111001) && ({row_reg, col_reg}<19'b0010100010100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100010100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100010100111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010100010100111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010100010101000000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010100010101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010100010101000010) && ({row_reg, col_reg}<19'b0010100010101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100010101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100010101001000) && ({row_reg, col_reg}<19'b0010100011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100011001010001) && ({row_reg, col_reg}<19'b0010100011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010100011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010100011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010100100000000000) && ({row_reg, col_reg}<19'b0010100100010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100100010110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010100100010110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100100010110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010100100010110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0010100100010111000) && ({row_reg, col_reg}<19'b0010100100010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100100010111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010100100010111101) && ({row_reg, col_reg}<19'b0010100100010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100100010111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100100011000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010100100011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010100100011000010) && ({row_reg, col_reg}<19'b0010100100011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100100011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100100011000110) && ({row_reg, col_reg}<19'b0010100100011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100100011010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010100100011010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010100100011011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100100011011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010100100011011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010100100011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010100100011011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010100100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100100011011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100100011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100100011100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0010100100011100001) && ({row_reg, col_reg}<19'b0010100100011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100100011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100100011100100) && ({row_reg, col_reg}<19'b0010100100011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100100011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100100011100111) && ({row_reg, col_reg}<19'b0010100100100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100100100100110) && ({row_reg, col_reg}<19'b0010100100100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100100100101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010100100100101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010100100100101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010100100100101100) && ({row_reg, col_reg}<19'b0010100100100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100100100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100100100111001) && ({row_reg, col_reg}<19'b0010100100100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100100100111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010100100100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0010100100100111111) && ({row_reg, col_reg}<19'b0010100100101000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100100101000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100100101000010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010100100101000011) && ({row_reg, col_reg}<19'b0010100101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100101001010001) && ({row_reg, col_reg}<19'b0010100101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010100101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010100101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010100110000000000) && ({row_reg, col_reg}<19'b0010100110010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100110010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100110010110010) && ({row_reg, col_reg}<19'b0010100110010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100110010110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010100110010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110010110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010100110010110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010100110010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100110010111001) && ({row_reg, col_reg}<19'b0010100110010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100110010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010100110010111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100110010111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110010111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010100110010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010100110011000000) && ({row_reg, col_reg}<19'b0010100110011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100110011000101) && ({row_reg, col_reg}<19'b0010100110011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100110011000111) && ({row_reg, col_reg}<19'b0010100110011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100110011010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100110011010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010100110011011000) && ({row_reg, col_reg}<19'b0010100110011011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110011011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010100110011011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100110011011100) && ({row_reg, col_reg}<19'b0010100110011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100110011011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100110011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110011100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100110011100001) && ({row_reg, col_reg}<19'b0010100110011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100110011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100110011100100) && ({row_reg, col_reg}<19'b0010100110011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100110011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010100110011100111) && ({row_reg, col_reg}<19'b0010100110100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100110100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010100110100100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010100110100101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0010100110100101001) && ({row_reg, col_reg}<19'b0010100110100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010100110100101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100110100101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010100110100101101) && ({row_reg, col_reg}<19'b0010100110100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010100110100111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010100110100111110) && ({row_reg, col_reg}<19'b0010100110101000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110101000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010100110101000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110101000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010100110101000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010100110101000100) && ({row_reg, col_reg}<19'b0010100111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010100111001010001) && ({row_reg, col_reg}<19'b0010100111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010100111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010100111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010101000000000000) && ({row_reg, col_reg}<19'b0010101000010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101000010110010) && ({row_reg, col_reg}<19'b0010101000010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000010110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101000010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000010110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101000010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101000010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101000010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101000010111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101000010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000010111101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101000010111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010101000010111111) && ({row_reg, col_reg}<19'b0010101000011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101000011000110) && ({row_reg, col_reg}<19'b0010101000011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101000011010011) && ({row_reg, col_reg}<19'b0010101000011010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101000011011000) && ({row_reg, col_reg}<19'b0010101000011011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000011011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000011011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010101000011011100) && ({row_reg, col_reg}<19'b0010101000011011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101000011011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101000011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000011100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010101000011100001) && ({row_reg, col_reg}<19'b0010101000011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101000011100100) && ({row_reg, col_reg}<19'b0010101000011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101000011100111) && ({row_reg, col_reg}<19'b0010101000100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101000100100001) && ({row_reg, col_reg}<19'b0010101000100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101000100100100) && ({row_reg, col_reg}<19'b0010101000100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000100100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101000100100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010101000100101000) && ({row_reg, col_reg}<19'b0010101000100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000100101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010101000100101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101000100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010101000100101110) && ({row_reg, col_reg}<19'b0010101000100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101000100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101000100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010101000100111110) && ({row_reg, col_reg}<19'b0010101000101000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000101000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000101000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101000101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000101000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101000101000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010101000101000101) && ({row_reg, col_reg}<19'b0010101001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010101001001010001) && ({row_reg, col_reg}<19'b0010101001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010101001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010101001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010101010000000000) && ({row_reg, col_reg}<19'b0010101010010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010010110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010101010010110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101010010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0010101010010110111) && ({row_reg, col_reg}<19'b0010101010010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010010111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010101010010111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010101010010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010010111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010101010010111110) && ({row_reg, col_reg}<19'b0010101010011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101010011010011) && ({row_reg, col_reg}<19'b0010101010011010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101010011011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101010011011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010011011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010101010011011011) && ({row_reg, col_reg}<19'b0010101010011011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010101010011011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101010011011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010011011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101010011100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010101010011100001) && ({row_reg, col_reg}<19'b0010101010011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101010011100100) && ({row_reg, col_reg}<19'b0010101010011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010011100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010101010011100111) && ({row_reg, col_reg}<19'b0010101010100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101010100100001) && ({row_reg, col_reg}<19'b0010101010100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101010100100100) && ({row_reg, col_reg}<19'b0010101010100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010101010100100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101010100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0010101010100101001) && ({row_reg, col_reg}<19'b0010101010100101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101010100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010100101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101010100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010101010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010101010100110000) && ({row_reg, col_reg}<19'b0010101010100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010101010100111011) && ({row_reg, col_reg}<19'b0010101010100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101010100111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101010100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010100111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101010101000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010101010101000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101010101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010101000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101010101000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101010101000110) && ({row_reg, col_reg}<19'b0010101011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010101011001010001) && ({row_reg, col_reg}<19'b0010101011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010101011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010101011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010101100000000000) && ({row_reg, col_reg}<19'b0010101100010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101100010110001) && ({row_reg, col_reg}<19'b0010101100010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100010110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010101100010110100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101100010110101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010101100010110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010101100010110111) && ({row_reg, col_reg}<19'b0010101100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101100010111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101100010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100010111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101100010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101100010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010101100011000000) && ({row_reg, col_reg}<19'b0010101100011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101100011010011) && ({row_reg, col_reg}<19'b0010101100011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100011011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010101100011011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101100011011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0010101100011011011) && ({row_reg, col_reg}<19'b0010101100011011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100011011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010101100011011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100011011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100011100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101100011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010101100011100010) && ({row_reg, col_reg}<19'b0010101100011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101100011100100) && ({row_reg, col_reg}<19'b0010101100011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100011100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010101100011100111) && ({row_reg, col_reg}<19'b0010101100100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100100100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010101100100100001) && ({row_reg, col_reg}<19'b0010101100100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101100100100100) && ({row_reg, col_reg}<19'b0010101100100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010101100100100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101100100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0010101100100101001) && ({row_reg, col_reg}<19'b0010101100100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010101100100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100100101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010101100100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101100100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100100101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010101100100110000) && ({row_reg, col_reg}<19'b0010101100100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101100100111001) && ({row_reg, col_reg}<19'b0010101100100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101100100111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101100100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100100111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0010101100101000000) && ({row_reg, col_reg}<19'b0010101100101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100101000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100101000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101100101000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010101100101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101100101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101100101001000) && ({row_reg, col_reg}<19'b0010101101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010101101001010001) && ({row_reg, col_reg}<19'b0010101101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010101101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010101101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010101110000000000) && ({row_reg, col_reg}<19'b0010101110010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101110010110001) && ({row_reg, col_reg}<19'b0010101110010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110010110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101110010110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010101110010110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101110010110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010101110010110111) && ({row_reg, col_reg}<19'b0010101110010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110010111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010101110010111010) && ({row_reg, col_reg}<19'b0010101110010111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010101110010111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010101110010111101) && ({row_reg, col_reg}<19'b0010101110010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110010111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010101110011000000) && ({row_reg, col_reg}<19'b0010101110011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010101110011010010) && ({row_reg, col_reg}<19'b0010101110011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101110011010100) && ({row_reg, col_reg}<19'b0010101110011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110011011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010101110011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101110011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010101110011011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101110011011101) && ({row_reg, col_reg}<19'b0010101110011011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101110011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101110011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101110011100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101110011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110011100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101110011100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010101110011100111) && ({row_reg, col_reg}<19'b0010101110100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110100100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010101110100100001) && ({row_reg, col_reg}<19'b0010101110100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101110100100100) && ({row_reg, col_reg}<19'b0010101110100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010101110100100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101110100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101110100101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010101110100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010101110100101011) && ({row_reg, col_reg}<19'b0010101110100101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101110100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010101110100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110100101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010101110100110000) && ({row_reg, col_reg}<19'b0010101110100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101110100111001) && ({row_reg, col_reg}<19'b0010101110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010101110100111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101110100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101110100111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101110101000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010101110101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110101000010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010101110101000011) && ({row_reg, col_reg}<19'b0010101110101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101110101000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010101110101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010101110101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010101110101001000) && ({row_reg, col_reg}<19'b0010101111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010101111001010001) && ({row_reg, col_reg}<19'b0010101111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010101111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010101111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010110000000000000) && ({row_reg, col_reg}<19'b0010110000010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010110000010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110000010110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010110000010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110000010110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110000010110110) && ({row_reg, col_reg}<19'b0010110000010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000010111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110000010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110000010111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110000010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110000010111101) && ({row_reg, col_reg}<19'b0010110000010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000011000000) && ({row_reg, col_reg}<19'b0010110000011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110000011111100) && ({row_reg, col_reg}<19'b0010110000011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000011111110) && ({row_reg, col_reg}<19'b0010110000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000100011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010110000100011001) && ({row_reg, col_reg}<19'b0010110000100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110000100011011) && ({row_reg, col_reg}<19'b0010110000100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000100011101) && ({row_reg, col_reg}<19'b0010110000100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000100011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110000100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000100100001) && ({row_reg, col_reg}<19'b0010110000100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110000100100100) && ({row_reg, col_reg}<19'b0010110000100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010110000100100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010110000100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010110000100101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110000100101010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010110000100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110000100101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010110000100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110000100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000100101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010110000100110000) && ({row_reg, col_reg}<19'b0010110000100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110000100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110000100111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010110000100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110000100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010110000101000000) && ({row_reg, col_reg}<19'b0010110000101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110000101000011) && ({row_reg, col_reg}<19'b0010110000101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110000101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110000101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000101000111) && ({row_reg, col_reg}<19'b0010110000101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110000101011110) && ({row_reg, col_reg}<19'b0010110000101100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000101100000) && ({row_reg, col_reg}<19'b0010110000101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110000101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000101101010) && ({row_reg, col_reg}<19'b0010110000101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000101101110) && ({row_reg, col_reg}<19'b0010110000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110000101111000) && ({row_reg, col_reg}<19'b0010110000101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000101111010) && ({row_reg, col_reg}<19'b0010110000110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110000110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000110000001) && ({row_reg, col_reg}<19'b0010110000110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110000110001000) && ({row_reg, col_reg}<19'b0010110000110001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110000110001101) && ({row_reg, col_reg}<19'b0010110001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110001001010001) && ({row_reg, col_reg}<19'b0010110001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010110001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010110001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010110010000000000) && ({row_reg, col_reg}<19'b0010110010010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010110010010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110010010110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010110010010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010010110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010110010010110110) && ({row_reg, col_reg}<19'b0010110010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010010111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110010010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010010111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110010010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110010010111101) && ({row_reg, col_reg}<19'b0010110010010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010011000000) && ({row_reg, col_reg}<19'b0010110010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010011111001) && ({row_reg, col_reg}<19'b0010110010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110010100011001) && ({row_reg, col_reg}<19'b0010110010100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110010100011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010100011101) && ({row_reg, col_reg}<19'b0010110010100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110010100011111) && ({row_reg, col_reg}<19'b0010110010100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010100100001) && ({row_reg, col_reg}<19'b0010110010100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010100100100) && ({row_reg, col_reg}<19'b0010110010100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010100100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110010100100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0010110010100101000) && ({row_reg, col_reg}<19'b0010110010100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010100101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010110010100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010100101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110010100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110010100110000) && ({row_reg, col_reg}<19'b0010110010100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010100111000) && ({row_reg, col_reg}<19'b0010110010100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010100111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110010100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010100111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010110010101000000) && ({row_reg, col_reg}<19'b0010110010101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110010101000011) && ({row_reg, col_reg}<19'b0010110010101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110010101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010101000111) && ({row_reg, col_reg}<19'b0010110010101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110010101100010) && ({row_reg, col_reg}<19'b0010110010101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010101100100) && ({row_reg, col_reg}<19'b0010110010101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110010101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110010101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110010101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010101101100) && ({row_reg, col_reg}<19'b0010110010101101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110010101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110010101101111) && ({row_reg, col_reg}<19'b0010110011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110011001010001) && ({row_reg, col_reg}<19'b0010110011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010110011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010110011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010110100000000000) && ({row_reg, col_reg}<19'b0010110100010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100010010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100010010001) && ({row_reg, col_reg}<19'b0010110100010010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100010011000) && ({row_reg, col_reg}<19'b0010110100010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010110100010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110100010110011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010110100010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110100010110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010110100010110110) && ({row_reg, col_reg}<19'b0010110100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100010111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110100010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110100010111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110100010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100010111101) && ({row_reg, col_reg}<19'b0010110100011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100100000000) && ({row_reg, col_reg}<19'b0010110100100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110100100011011) && ({row_reg, col_reg}<19'b0010110100100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100100011101) && ({row_reg, col_reg}<19'b0010110100100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100100100001) && ({row_reg, col_reg}<19'b0010110100100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110100100100011) && ({row_reg, col_reg}<19'b0010110100100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110100100100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010110100100101000) && ({row_reg, col_reg}<19'b0010110100100101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010110100100101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110100100101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110100100101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010110100100101101) && ({row_reg, col_reg}<19'b0010110100100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100100110000) && ({row_reg, col_reg}<19'b0010110100100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110100100110100) && ({row_reg, col_reg}<19'b0010110100100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110100100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110100100111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110100100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110100100111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010110100101000000) && ({row_reg, col_reg}<19'b0010110100101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110100101000011) && ({row_reg, col_reg}<19'b0010110100101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110100101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110100101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100101000111) && ({row_reg, col_reg}<19'b0010110100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110100101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100101100100) && ({row_reg, col_reg}<19'b0010110100101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110100101101100) && ({row_reg, col_reg}<19'b0010110100101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100101101110) && ({row_reg, col_reg}<19'b0010110100110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110100110001110) && ({row_reg, col_reg}<19'b0010110100110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110100110010000) && ({row_reg, col_reg}<19'b0010110101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110101001010001) && ({row_reg, col_reg}<19'b0010110101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010110101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010110101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010110110000000000) && ({row_reg, col_reg}<19'b0010110110010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110110010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110010110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010110110010110011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010110110010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110110010110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010110110010110110) && ({row_reg, col_reg}<19'b0010110110010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110110010111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110110010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110110010111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110110010111100) && ({row_reg, col_reg}<19'b0010110110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110110011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110110100000000) && ({row_reg, col_reg}<19'b0010110110100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110110100100001) && ({row_reg, col_reg}<19'b0010110110100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110110100100011) && ({row_reg, col_reg}<19'b0010110110100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110110100100101) && ({row_reg, col_reg}<19'b0010110110100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110100100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110110100101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010110110100101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110110100101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010110110100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010110110100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110110100101101) && ({row_reg, col_reg}<19'b0010110110100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110110100101111) && ({row_reg, col_reg}<19'b0010110110100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110110100110110) && ({row_reg, col_reg}<19'b0010110110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110110100111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110110100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110110100111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010110110101000000) && ({row_reg, col_reg}<19'b0010110110101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110110101000011) && ({row_reg, col_reg}<19'b0010110110101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110110101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010110110101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110110101000111) && ({row_reg, col_reg}<19'b0010110110101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110110101011011) && ({row_reg, col_reg}<19'b0010110110101100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110110101100000) && ({row_reg, col_reg}<19'b0010110110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010110110101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110110101111001) && ({row_reg, col_reg}<19'b0010110110110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110110110001000) && ({row_reg, col_reg}<19'b0010110110110001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010110110110001010) && ({row_reg, col_reg}<19'b0010110110110001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010110110110001101) && ({row_reg, col_reg}<19'b0010110111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010110111001010001) && ({row_reg, col_reg}<19'b0010110111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010110111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010110111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010111000000000000) && ({row_reg, col_reg}<19'b0010111000010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111000010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000010110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111000010110011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010111000010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111000010110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010111000010110110) && ({row_reg, col_reg}<19'b0010111000010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111000010111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111000010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111000010111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010111000010111100) && ({row_reg, col_reg}<19'b0010111000010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000010111111) && ({row_reg, col_reg}<19'b0010111000100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000100100001) && ({row_reg, col_reg}<19'b0010111000100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111000100100100) && ({row_reg, col_reg}<19'b0010111000100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000100100110) && ({row_reg, col_reg}<19'b0010111000100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111000100101001) && ({row_reg, col_reg}<19'b0010111000100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111000100101011) && ({row_reg, col_reg}<19'b0010111000100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111000100101101) && ({row_reg, col_reg}<19'b0010111000100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000100101111) && ({row_reg, col_reg}<19'b0010111000100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111000100110100) && ({row_reg, col_reg}<19'b0010111000100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000100110110) && ({row_reg, col_reg}<19'b0010111000100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000100111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111000100111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111000100111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010111000100111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010111000101000000) && ({row_reg, col_reg}<19'b0010111000101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111000101000011) && ({row_reg, col_reg}<19'b0010111000101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111000101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111000101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000101000111) && ({row_reg, col_reg}<19'b0010111000101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111000101100000) && ({row_reg, col_reg}<19'b0010111000101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000101100010) && ({row_reg, col_reg}<19'b0010111000101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111000101100110) && ({row_reg, col_reg}<19'b0010111000101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111000101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111000101101001) && ({row_reg, col_reg}<19'b0010111000101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000101101011) && ({row_reg, col_reg}<19'b0010111000101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111000101101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111000101110000) && ({row_reg, col_reg}<19'b0010111000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000101111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111000101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000101111010) && ({row_reg, col_reg}<19'b0010111000110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111000110000000) && ({row_reg, col_reg}<19'b0010111000110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000110000010) && ({row_reg, col_reg}<19'b0010111000110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111000110001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000110001011) && ({row_reg, col_reg}<19'b0010111000110001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111000110001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111000110001110) && ({row_reg, col_reg}<19'b0010111001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111001001010001) && ({row_reg, col_reg}<19'b0010111001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010111001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010111001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010111010000000000) && ({row_reg, col_reg}<19'b0010111010010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111010010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010010110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010111010010110011) && ({row_reg, col_reg}<19'b0010111010010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111010010110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010111010010110110) && ({row_reg, col_reg}<19'b0010111010010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111010010111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010111010010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111010010111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010111010010111100) && ({row_reg, col_reg}<19'b0010111010010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111010010111111) && ({row_reg, col_reg}<19'b0010111010100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010100011010) && ({row_reg, col_reg}<19'b0010111010100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111010100011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010111010100011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111010100011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010100100000) && ({row_reg, col_reg}<19'b0010111010100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111010100100100) && ({row_reg, col_reg}<19'b0010111010100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010100100110) && ({row_reg, col_reg}<19'b0010111010100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111010100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111010100101011) && ({row_reg, col_reg}<19'b0010111010100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010100101110) && ({row_reg, col_reg}<19'b0010111010100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010100110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010111010100110101) && ({row_reg, col_reg}<19'b0010111010100110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010111010100110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111010100111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010111010100111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010111010100111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010111010100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111010100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0010111010100111101) && ({row_reg, col_reg}<19'b0010111010100111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111010100111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0010111010101000000) && ({row_reg, col_reg}<19'b0010111010101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111010101000011) && ({row_reg, col_reg}<19'b0010111010101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111010101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111010101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010101000111) && ({row_reg, col_reg}<19'b0010111010101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111010101011000) && ({row_reg, col_reg}<19'b0010111010101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010101011010) && ({row_reg, col_reg}<19'b0010111010101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010101100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010101100001) && ({row_reg, col_reg}<19'b0010111010101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111010101101000) && ({row_reg, col_reg}<19'b0010111010101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010101101011) && ({row_reg, col_reg}<19'b0010111010101101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010101110000) && ({row_reg, col_reg}<19'b0010111010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010101111001) && ({row_reg, col_reg}<19'b0010111010101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111010101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010101111100) && ({row_reg, col_reg}<19'b0010111010101111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111010101111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111010101111111) && ({row_reg, col_reg}<19'b0010111010110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111010110001100) && ({row_reg, col_reg}<19'b0010111010110001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111010110001110) && ({row_reg, col_reg}<19'b0010111011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111011001010001) && ({row_reg, col_reg}<19'b0010111011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010111011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010111011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010111100000000000) && ({row_reg, col_reg}<19'b0010111100010010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100010010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111100010010011) && ({row_reg, col_reg}<19'b0010111100010010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111100010010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111100010010110) && ({row_reg, col_reg}<19'b0010111100010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111100010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100010110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010111100010110011) && ({row_reg, col_reg}<19'b0010111100010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111100010110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010111100010110110) && ({row_reg, col_reg}<19'b0010111100010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100010111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111100010111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010111100010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111100010111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010111100010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111100010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111100010111111) && ({row_reg, col_reg}<19'b0010111100011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100011111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111100011111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100011111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111100011111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010111100011111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010111100100000000) && ({row_reg, col_reg}<19'b0010111100100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100100011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010111100100011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111100100011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111100100011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111100100011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111100100011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010111100100011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111100100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111100100100001) && ({row_reg, col_reg}<19'b0010111100100100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111100100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111100100100101) && ({row_reg, col_reg}<19'b0010111100100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111100100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111100100101000) && ({row_reg, col_reg}<19'b0010111100100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111100100101011) && ({row_reg, col_reg}<19'b0010111100100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111100100101110) && ({row_reg, col_reg}<19'b0010111100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100100110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111100100110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100100110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111100100110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111100100110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111100100111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010111100100111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0010111100100111010) && ({row_reg, col_reg}<19'b0010111100100111101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010111100100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111100100111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010111100100111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010111100101000000) && ({row_reg, col_reg}<19'b0010111100101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111100101000011) && ({row_reg, col_reg}<19'b0010111100101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111100101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111100101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111100101000111) && ({row_reg, col_reg}<19'b0010111100101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111100101011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111100101011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010111100101011111) && ({row_reg, col_reg}<19'b0010111100101100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010111100101100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010111100101100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010111100101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111100101100110) && ({row_reg, col_reg}<19'b0010111100101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111100101101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111100101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111100101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111100101101101) && ({row_reg, col_reg}<19'b0010111100101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100101111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111100101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100101111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111100101111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111100101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100101111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010111100110000000) && ({row_reg, col_reg}<19'b0010111100110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100110000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111100110000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010111100110000100) && ({row_reg, col_reg}<19'b0010111100110000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010111100110000110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010111100110000111) && ({row_reg, col_reg}<19'b0010111100110001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010111100110001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111100110001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111100110001011) && ({row_reg, col_reg}<19'b0010111100110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111100110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111100110010000) && ({row_reg, col_reg}<19'b0010111101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111101001010001) && ({row_reg, col_reg}<19'b0010111101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010111101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010111101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0010111110000000000) && ({row_reg, col_reg}<19'b0010111110010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110010010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111110010010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0010111110010010011) && ({row_reg, col_reg}<19'b0010111110010010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010111110010010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111110010010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111110010010111) && ({row_reg, col_reg}<19'b0010111110010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111110010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110010110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0010111110010110011) && ({row_reg, col_reg}<19'b0010111110010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110010110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0010111110010110110) && ({row_reg, col_reg}<19'b0010111110010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110010111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111110010111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010111110010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110010111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010111110010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111110010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111110010111111) && ({row_reg, col_reg}<19'b0010111110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111110011111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110011111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010111110011111101) && ({row_reg, col_reg}<19'b0010111110011111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110011111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010111110100000000) && ({row_reg, col_reg}<19'b0010111110100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110100011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110100011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010111110100011011) && ({row_reg, col_reg}<19'b0010111110100011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111110100011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111110100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111110100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111110100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111110100100100) && ({row_reg, col_reg}<19'b0010111110100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111110100100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111110100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111110100101001) && ({row_reg, col_reg}<19'b0010111110100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111110100110000) && ({row_reg, col_reg}<19'b0010111110100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111110100110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010111110100110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0010111110100110101) && ({row_reg, col_reg}<19'b0010111110100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110100111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010111110100111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110100111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010111110100111100) && ({row_reg, col_reg}<19'b0010111110100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111110100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0010111110100111111) && ({row_reg, col_reg}<19'b0010111110101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0010111110101000011) && ({row_reg, col_reg}<19'b0010111110101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111110101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111110101000111) && ({row_reg, col_reg}<19'b0010111110101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0010111110101011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010111110101011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111110101011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010111110101011111) && ({row_reg, col_reg}<19'b0010111110101100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110101100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010111110101100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111110101100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010111110101100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0010111110101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111110101101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0010111110101101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111110101101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111110101101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110101101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0010111110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111110101101111) && ({row_reg, col_reg}<19'b0010111110101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110101111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111110101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110101111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0010111110101111100) && ({row_reg, col_reg}<19'b0010111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110101111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111110101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110110000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0010111110110000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010111110110000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0010111110110000011) && ({row_reg, col_reg}<19'b0010111110110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110110000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0010111110110001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0010111110110001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111110110001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0010111110110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111110110001100) && ({row_reg, col_reg}<19'b0010111110110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0010111110110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0010111110110010000) && ({row_reg, col_reg}<19'b0010111111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0010111111001010001) && ({row_reg, col_reg}<19'b0010111111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0010111111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0010111111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011000000000000000) && ({row_reg, col_reg}<19'b0011000000010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000010010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000000010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011000000010010011) && ({row_reg, col_reg}<19'b0011000000010010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000010010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000010010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000010010111) && ({row_reg, col_reg}<19'b0011000000010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000000010110011) && ({row_reg, col_reg}<19'b0011000000010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000000010110110) && ({row_reg, col_reg}<19'b0011000000010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000000010111001) && ({row_reg, col_reg}<19'b0011000000010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000010111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000000010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000010111101) && ({row_reg, col_reg}<19'b0011000000010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000011000000) && ({row_reg, col_reg}<19'b0011000000011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000011010011) && ({row_reg, col_reg}<19'b0011000000011010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000011010110) && ({row_reg, col_reg}<19'b0011000000011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000000011011110) && ({row_reg, col_reg}<19'b0011000000011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000011100001) && ({row_reg, col_reg}<19'b0011000000011100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000000011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000000011100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000000011100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000011100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000000011100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000000011101000) && ({row_reg, col_reg}<19'b0011000000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000000011101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000000011101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000000011101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000011101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000000011101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000000011110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000000011110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000011110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011000000011110011) && ({row_reg, col_reg}<19'b0011000000011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000011110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000011110111) && ({row_reg, col_reg}<19'b0011000000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000011111010) && ({row_reg, col_reg}<19'b0011000000011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000011111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000011111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000000011111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000011111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000100000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000000100000010) && ({row_reg, col_reg}<19'b0011000000100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000100000101) && ({row_reg, col_reg}<19'b0011000000100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100000111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000000100001000) && ({row_reg, col_reg}<19'b0011000000100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000100010011) && ({row_reg, col_reg}<19'b0011000000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000000100011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000000100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000100011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000100011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000000100011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000100011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000100011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011000000100100000) && ({row_reg, col_reg}<19'b0011000000100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000100100100) && ({row_reg, col_reg}<19'b0011000000100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000000100101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000100101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000000100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000000100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000000100110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000000100110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000100110101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000100110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011000000100110111) && ({row_reg, col_reg}<19'b0011000000100111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000000100111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000000100111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000000100111100) && ({row_reg, col_reg}<19'b0011000000100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000000100111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011000000101000000) && ({row_reg, col_reg}<19'b0011000000101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000000101000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011000000101000100) && ({row_reg, col_reg}<19'b0011000000101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000101000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000000101000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000101001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000101001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000000101001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000000101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000000101001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000101001101) && ({row_reg, col_reg}<19'b0011000000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000101001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000000101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000101010001) && ({row_reg, col_reg}<19'b0011000000101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000000101010011) && ({row_reg, col_reg}<19'b0011000000101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000000101010101) && ({row_reg, col_reg}<19'b0011000000101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000000101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000000101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000000101011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011000000101011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011000000101011101) && ({row_reg, col_reg}<19'b0011000000101011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011000000101011111) && ({row_reg, col_reg}<19'b0011000000101100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000000101100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011000000101100011) && ({row_reg, col_reg}<19'b0011000000101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000101100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000101100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000000101101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011000000101101001) && ({row_reg, col_reg}<19'b0011000000101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000101101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000000101101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000101101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000000101101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011000000101101111) && ({row_reg, col_reg}<19'b0011000000101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000000101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000101111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000000101111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000101111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000000101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000110000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000110000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000000110000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000000110000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000000110000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000110000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000110000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000110000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000000110001000) && ({row_reg, col_reg}<19'b0011000000110001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000110001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000110001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000000110001101) && ({row_reg, col_reg}<19'b0011000000110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000000110001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000000110010000) && ({row_reg, col_reg}<19'b0011000001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000001001010001) && ({row_reg, col_reg}<19'b0011000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011000001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011000001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011000010000000000) && ({row_reg, col_reg}<19'b0011000010010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010010010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000010010010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000010010010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000010010010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000010010010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000010010010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010010010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000010010010111) && ({row_reg, col_reg}<19'b0011000010010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000010010110011) && ({row_reg, col_reg}<19'b0011000010010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000010010110110) && ({row_reg, col_reg}<19'b0011000010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000010010111001) && ({row_reg, col_reg}<19'b0011000010010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010010111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000010010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000010010111101) && ({row_reg, col_reg}<19'b0011000010010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010011000000) && ({row_reg, col_reg}<19'b0011000010011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010011010011) && ({row_reg, col_reg}<19'b0011000010011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010011011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000010011011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011000010011011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010011011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000010011011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000010011011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011000010011011111) && ({row_reg, col_reg}<19'b0011000010011100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000010011100001) && ({row_reg, col_reg}<19'b0011000010011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011000010011100011) && ({row_reg, col_reg}<19'b0011000010011100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011000010011100101) && ({row_reg, col_reg}<19'b0011000010011101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010011101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011000010011101101) && ({row_reg, col_reg}<19'b0011000010011101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000010011101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000010011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010011110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000010011110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000010011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000010011110101) && ({row_reg, col_reg}<19'b0011000010011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010011110111) && ({row_reg, col_reg}<19'b0011000010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010011111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000010011111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000010011111100) && ({row_reg, col_reg}<19'b0011000010011111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000010011111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011000010011111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000010100000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000010100000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000010100000010) && ({row_reg, col_reg}<19'b0011000010100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010100000101) && ({row_reg, col_reg}<19'b0011000010100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000010100001000) && ({row_reg, col_reg}<19'b0011000010100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010100010011) && ({row_reg, col_reg}<19'b0011000010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010100011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011000010100011001) && ({row_reg, col_reg}<19'b0011000010100011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000010100011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000010100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010100011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000010100011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010100011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011000010100100000) && ({row_reg, col_reg}<19'b0011000010100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000010100100111) && ({row_reg, col_reg}<19'b0011000010100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000010100101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010100101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011000010100101011) && ({row_reg, col_reg}<19'b0011000010100101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000010100101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000010100101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011000010100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000010100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000010100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010100110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000010100110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000010100110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000010100110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000010100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010100110111) && ({row_reg, col_reg}<19'b0011000010100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000010100111001) && ({row_reg, col_reg}<19'b0011000010100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000010100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000010100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010100111101) && ({row_reg, col_reg}<19'b0011000010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010101000001) && ({row_reg, col_reg}<19'b0011000010101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010101000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011000010101000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000010101000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000010101000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011000010101000111) && ({row_reg, col_reg}<19'b0011000010101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010101001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000010101001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000010101001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011000010101001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010101001111) && ({row_reg, col_reg}<19'b0011000010101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000010101010011) && ({row_reg, col_reg}<19'b0011000010101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010101010101) && ({row_reg, col_reg}<19'b0011000010101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000010101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010101011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000010101011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011000010101011011) && ({row_reg, col_reg}<19'b0011000010101011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010101011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000010101011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010101011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000010101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010101100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000010101100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000010101100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000010101100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010101100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000010101100110) && ({row_reg, col_reg}<19'b0011000010101101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010101101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000010101101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011000010101101100) && ({row_reg, col_reg}<19'b0011000010101101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010101101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000010101101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000010101110000) && ({row_reg, col_reg}<19'b0011000010101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000010101111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000010101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010101111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000010101111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011000010101111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011000010101111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000010101111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000010110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010110000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000010110000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000010110000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011000010110000100) && ({row_reg, col_reg}<19'b0011000010110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000010110000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000010110000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011000010110001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000010110001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011000010110001010) && ({row_reg, col_reg}<19'b0011000010110001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000010110001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000010110001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011000010110001110) && ({row_reg, col_reg}<19'b0011000010110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000010110010000) && ({row_reg, col_reg}<19'b0011000011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000011001010001) && ({row_reg, col_reg}<19'b0011000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011000011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011000011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011000100000000000) && ({row_reg, col_reg}<19'b0011000100010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100010010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000100010010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011000100010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000100010010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100010010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000100010010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011000100010010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000100010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000100010011000) && ({row_reg, col_reg}<19'b0011000100010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000100010110011) && ({row_reg, col_reg}<19'b0011000100010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000100010110110) && ({row_reg, col_reg}<19'b0011000100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100010111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000100010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100010111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011000100010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000100010111101) && ({row_reg, col_reg}<19'b0011000100010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000100011000000) && ({row_reg, col_reg}<19'b0011000100011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100011011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000100011011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100011011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011000100011011011) && ({row_reg, col_reg}<19'b0011000100011100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100011100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011000100011100001) && ({row_reg, col_reg}<19'b0011000100011100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100011100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000100011100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100011101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011000100011101001) && ({row_reg, col_reg}<19'b0011000100011101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000100011101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000100011101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000100011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011000100011110001) && ({row_reg, col_reg}<19'b0011000100011110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100011110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000100011110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000100011110101) && ({row_reg, col_reg}<19'b0011000100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100011111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000100011111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000100011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100011111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000100011111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000100100000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000100100000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011000100100000010) && ({row_reg, col_reg}<19'b0011000100100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000100100000101) && ({row_reg, col_reg}<19'b0011000100100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000100100001000) && ({row_reg, col_reg}<19'b0011000100100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000100100010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000100100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000100100011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000100100011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000100100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000100100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100100011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100100011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000100100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000100100100001) && ({row_reg, col_reg}<19'b0011000100100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000100100101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000100100101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100100101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000100100101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000100100101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000100100101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000100100101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000100100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000100100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100100110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011000100100110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100100110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000100100110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000100100110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000100100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000100100111000) && ({row_reg, col_reg}<19'b0011000100100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000100100111101) && ({row_reg, col_reg}<19'b0011000100100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000100101000001) && ({row_reg, col_reg}<19'b0011000100101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000100101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000100101000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000100101000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000100101000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000100101001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000100101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100101001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000100101001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000100101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100101001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000100101001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011000100101001111) && ({row_reg, col_reg}<19'b0011000100101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000100101010011) && ({row_reg, col_reg}<19'b0011000100101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000100101010101) && ({row_reg, col_reg}<19'b0011000100101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000100101010111) && ({row_reg, col_reg}<19'b0011000100101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000100101011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011000100101011010) && ({row_reg, col_reg}<19'b0011000100101011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100101011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100101011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011000100101011110) && ({row_reg, col_reg}<19'b0011000100101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000100101100001) && ({row_reg, col_reg}<19'b0011000100101100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000100101100011) && ({row_reg, col_reg}<19'b0011000100101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100101100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000100101100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011000100101100111) && ({row_reg, col_reg}<19'b0011000100101101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100101101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000100101101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000100101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000100101101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000100101101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100101101110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100101101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000100101110000) && ({row_reg, col_reg}<19'b0011000100101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100101111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000100101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100101111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011000100101111100) && ({row_reg, col_reg}<19'b0011000100101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100101111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011000100101111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000100110000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100110000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100110000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000100110000011) && ({row_reg, col_reg}<19'b0011000100110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000100110000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000100110001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000100110001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000100110001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100110001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100110001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100110001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000100110001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011000100110001111) && ({row_reg, col_reg}<19'b0011000101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000101001010001) && ({row_reg, col_reg}<19'b0011000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011000101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011000101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011000110000000000) && ({row_reg, col_reg}<19'b0011000110010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110010010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110010010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011000110010010010) && ({row_reg, col_reg}<19'b0011000110010010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000110010010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110010010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000110010010110) && ({row_reg, col_reg}<19'b0011000110010011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110010011000) && ({row_reg, col_reg}<19'b0011000110010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000110010110011) && ({row_reg, col_reg}<19'b0011000110010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000110010110110) && ({row_reg, col_reg}<19'b0011000110010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110010111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000110010111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000110010111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000110010111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000110010111101) && ({row_reg, col_reg}<19'b0011000110010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110011000000) && ({row_reg, col_reg}<19'b0011000110011010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110011010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000110011011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000110011011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000110011011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110011011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000110011011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000110011011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000110011011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000110011011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000110011100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011000110011100001) && ({row_reg, col_reg}<19'b0011000110011100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011000110011100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011000110011100100) && ({row_reg, col_reg}<19'b0011000110011100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000110011100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000110011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110011101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000110011101001) && ({row_reg, col_reg}<19'b0011000110011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110011110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000110011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110011110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000110011110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000110011110101) && ({row_reg, col_reg}<19'b0011000110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110011111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110011111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000110011111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000110011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110011111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000110100000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110100000011) && ({row_reg, col_reg}<19'b0011000110100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110100010100) && ({row_reg, col_reg}<19'b0011000110100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000110100010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011000110100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110100011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000110100011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011000110100011011) && ({row_reg, col_reg}<19'b0011000110100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110100011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011000110100011110) && ({row_reg, col_reg}<19'b0011000110100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110100100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011000110100100001) && ({row_reg, col_reg}<19'b0011000110100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110100101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011000110100101001) && ({row_reg, col_reg}<19'b0011000110100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110100101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000110100101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000110100101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000110100101110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000110100101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011000110100110000) && ({row_reg, col_reg}<19'b0011000110100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110100110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000110100110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011000110100110100) && ({row_reg, col_reg}<19'b0011000110100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110100110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000110100110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011000110100111000) && ({row_reg, col_reg}<19'b0011000110100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110100111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000110100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011000110100111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000110101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110101000001) && ({row_reg, col_reg}<19'b0011000110101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110101001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110101001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011000110101001100) && ({row_reg, col_reg}<19'b0011000110101001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011000110101001111) && ({row_reg, col_reg}<19'b0011000110101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110101010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110101010100) && ({row_reg, col_reg}<19'b0011000110101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110101010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000110101011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000110101011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000110101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110101011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000110101011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000110101011101) && ({row_reg, col_reg}<19'b0011000110101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011000110101100000) && ({row_reg, col_reg}<19'b0011000110101100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000110101100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000110101100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011000110101100100) && ({row_reg, col_reg}<19'b0011000110101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110101100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011000110101100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011000110101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110101101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000110101101010) && ({row_reg, col_reg}<19'b0011000110101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110101101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000110101101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011000110101101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110101101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011000110101110000) && ({row_reg, col_reg}<19'b0011000110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110101111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000110101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011000110101111100) && ({row_reg, col_reg}<19'b0011000110101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110101111111) && ({row_reg, col_reg}<19'b0011000110110000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011000110110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110110000010) && ({row_reg, col_reg}<19'b0011000110110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110110000110) && ({row_reg, col_reg}<19'b0011000110110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110110001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011000110110001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011000110110001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011000110110001100) && ({row_reg, col_reg}<19'b0011000110110001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110110001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000110110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011000110110010000) && ({row_reg, col_reg}<19'b0011000111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011000111001010001) && ({row_reg, col_reg}<19'b0011000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011000111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011000111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011001000000000000) && ({row_reg, col_reg}<19'b0011001000010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000010010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011001000010010010) && ({row_reg, col_reg}<19'b0011001000010010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001000010010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011001000010010101) && ({row_reg, col_reg}<19'b0011001000010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001000010110011) && ({row_reg, col_reg}<19'b0011001000010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001000010110110) && ({row_reg, col_reg}<19'b0011001000010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000010111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000010111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001000010111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001000010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011001000010111101) && ({row_reg, col_reg}<19'b0011001000011010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000011010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000011010100) && ({row_reg, col_reg}<19'b0011001000011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000011010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001000011010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001000011011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000011011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001000011011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001000011011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001000011011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001000011011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000011011110) && ({row_reg, col_reg}<19'b0011001000011101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000011101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000011101001) && ({row_reg, col_reg}<19'b0011001000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001000011110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001000011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000011110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001000011110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001000011110101) && ({row_reg, col_reg}<19'b0011001000011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001000011111010) && ({row_reg, col_reg}<19'b0011001000011111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001000011111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001000011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001000011111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001000100000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000100000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001000100000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001000100000011) && ({row_reg, col_reg}<19'b0011001000100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000100010100) && ({row_reg, col_reg}<19'b0011001000100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000100010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001000100010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001000100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000100011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000100011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011001000100011011) && ({row_reg, col_reg}<19'b0011001000100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000100011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001000100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001000100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000100100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001000100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000100100010) && ({row_reg, col_reg}<19'b0011001000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001000100101001) && ({row_reg, col_reg}<19'b0011001000100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001000100101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001000100101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001000100101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001000100101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001000100110000) && ({row_reg, col_reg}<19'b0011001000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001000100110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001000100110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001000100110101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001000100110110) && ({row_reg, col_reg}<19'b0011001000100111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000100111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001000100111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001000100111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001000100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001000101000001) && ({row_reg, col_reg}<19'b0011001000101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000101000100) && ({row_reg, col_reg}<19'b0011001000101000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011001000101000110) && ({row_reg, col_reg}<19'b0011001000101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001000101001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001000101001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001000101001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001000101001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001000101001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001000101001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001000101001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001000101001111) && ({row_reg, col_reg}<19'b0011001000101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000101010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000101010100) && ({row_reg, col_reg}<19'b0011001000101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001000101010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000101011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000101011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001000101011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001000101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000101011100) && ({row_reg, col_reg}<19'b0011001000101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000101011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001000101011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001000101100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000101100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001000101100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001000101100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000101100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001000101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000101100111) && ({row_reg, col_reg}<19'b0011001000101101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001000101101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001000101101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001000101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000101101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001000101101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001000101101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000101101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001000101110000) && ({row_reg, col_reg}<19'b0011001000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000101111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001000101111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001000101111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001000101111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001000101111100) && ({row_reg, col_reg}<19'b0011001000101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001000101111111) && ({row_reg, col_reg}<19'b0011001000110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000110000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001000110000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001000110000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001000110000111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001000110001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001000110001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001000110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001000110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001000110001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001000110001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000110001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001000110001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001000110010000) && ({row_reg, col_reg}<19'b0011001001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001001001010001) && ({row_reg, col_reg}<19'b0011001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011001001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011001001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011001010000000000) && ({row_reg, col_reg}<19'b0011001010010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010010010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001010010010010) && ({row_reg, col_reg}<19'b0011001010010010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001010010010100) && ({row_reg, col_reg}<19'b0011001010010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001010010110011) && ({row_reg, col_reg}<19'b0011001010010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001010010110110) && ({row_reg, col_reg}<19'b0011001010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001010010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001010010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010010111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011001010010111101) && ({row_reg, col_reg}<19'b0011001010011010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010011010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001010011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010011010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010011010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001010011010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001010011011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010011011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001010011011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001010011011011) && ({row_reg, col_reg}<19'b0011001010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001010011011101) && ({row_reg, col_reg}<19'b0011001010011011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001010011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010011100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010011100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001010011100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001010011100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001010011100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001010011100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001010011101000) && ({row_reg, col_reg}<19'b0011001010011101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010011101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010011101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001010011101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001010011101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010011101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001010011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011001010011110001) && ({row_reg, col_reg}<19'b0011001010011110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010011110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001010011110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001010011110101) && ({row_reg, col_reg}<19'b0011001010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010011111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001010011111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001010011111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010011111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001010100000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010100000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001010100000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011001010100000011) && ({row_reg, col_reg}<19'b0011001010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001010100010001) && ({row_reg, col_reg}<19'b0011001010100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001010100010100) && ({row_reg, col_reg}<19'b0011001010100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010100010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010100010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001010100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001010100011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001010100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010100100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001010100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001010100100010) && ({row_reg, col_reg}<19'b0011001010100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001010100101001) && ({row_reg, col_reg}<19'b0011001010100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010100101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001010100101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001010100101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001010100101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001010100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001010100110001) && ({row_reg, col_reg}<19'b0011001010100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010100110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001010100110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001010100110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001010100110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001010100111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001010100111010) && ({row_reg, col_reg}<19'b0011001010100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010100111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001010100111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001010100111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001010101000001) && ({row_reg, col_reg}<19'b0011001010101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010101000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010101000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001010101000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001010101000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001010101000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011001010101001000) && ({row_reg, col_reg}<19'b0011001010101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001010101001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010101001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011001010101001111) && ({row_reg, col_reg}<19'b0011001010101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010101010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010101010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001010101011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010101011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001010101011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001010101011011) && ({row_reg, col_reg}<19'b0011001010101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010101011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001010101011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001010101011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001010101100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001010101100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010101100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011001010101100011) && ({row_reg, col_reg}<19'b0011001010101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010101100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001010101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010101100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010101101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010101101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001010101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010101101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001010101101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010101101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011001010101110000) && ({row_reg, col_reg}<19'b0011001010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010101111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001010101111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001010101111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001010101111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010101111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001010101111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001010101111111) && ({row_reg, col_reg}<19'b0011001010110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001010110000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001010110000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001010110000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001010110000110) && ({row_reg, col_reg}<19'b0011001010110001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010110001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001010110001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001010110001010) && ({row_reg, col_reg}<19'b0011001010110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001010110001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001010110001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001010110001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010110001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011001010110010000) && ({row_reg, col_reg}<19'b0011001011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001011001010001) && ({row_reg, col_reg}<19'b0011001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011001011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011001011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011001100000000000) && ({row_reg, col_reg}<19'b0011001100010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001100010110011) && ({row_reg, col_reg}<19'b0011001100010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001100010110110) && ({row_reg, col_reg}<19'b0011001100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001100010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001100010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100010111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001100010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001100010111111) && ({row_reg, col_reg}<19'b0011001100011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001100011010001) && ({row_reg, col_reg}<19'b0011001100011010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100011010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001100011010100) && ({row_reg, col_reg}<19'b0011001100011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100011010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001100011010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001100011011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001100011011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100011011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001100011011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100011011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011001100011011110) && ({row_reg, col_reg}<19'b0011001100011100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100011100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011001100011100001) && ({row_reg, col_reg}<19'b0011001100011100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100011100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001100011100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001100011100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011001100011100110) && ({row_reg, col_reg}<19'b0011001100011101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100011101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001100011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100011101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100011101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001100011101110) && ({row_reg, col_reg}<19'b0011001100011110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100011110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001100011110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001100011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001100011110101) && ({row_reg, col_reg}<19'b0011001100011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001100011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001100011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100011111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001100011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100011111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001100011111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100011111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001100100000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100100000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001100100000010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011001100100000011) && ({row_reg, col_reg}<19'b0011001100100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001100100000101) && ({row_reg, col_reg}<19'b0011001100100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001100100000111) && ({row_reg, col_reg}<19'b0011001100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001100100010001) && ({row_reg, col_reg}<19'b0011001100100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001100100010100) && ({row_reg, col_reg}<19'b0011001100100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100100010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001100100010111) && ({row_reg, col_reg}<19'b0011001100100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100100011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001100100011010) && ({row_reg, col_reg}<19'b0011001100100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001100100011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100100100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001100100100010) && ({row_reg, col_reg}<19'b0011001100100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100100101010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001100100101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001100100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001100100101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001100100101110) && ({row_reg, col_reg}<19'b0011001100100110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011001100100110000) && ({row_reg, col_reg}<19'b0011001100100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001100100110010) && ({row_reg, col_reg}<19'b0011001100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100100111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001100100111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001100100111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001100100111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001100100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001100100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001100101000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001100101000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011001100101000100) && ({row_reg, col_reg}<19'b0011001100101000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011001100101000110) && ({row_reg, col_reg}<19'b0011001100101001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100101001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001100101001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100101001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001100101001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001100101001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001100101001111) && ({row_reg, col_reg}<19'b0011001100101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001100101010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001100101010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100101011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001100101011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011001100101011010) && ({row_reg, col_reg}<19'b0011001100101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100101011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001100101011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001100101011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001100101011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001100101100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011001100101100001) && ({row_reg, col_reg}<19'b0011001100101100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001100101100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001100101100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001100101100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100101100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001100101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001100101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001100101101010) && ({row_reg, col_reg}<19'b0011001100101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001100101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100101101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001100101101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011001100101101111) && ({row_reg, col_reg}<19'b0011001100101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100101111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001100101111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001100101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100101111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001100101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001100101111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001100101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001100110000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001100110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001100110000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001100110000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011001100110000101) && ({row_reg, col_reg}<19'b0011001100110001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100110001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001100110001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001100110001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001100110001011) && ({row_reg, col_reg}<19'b0011001100110001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001100110001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001100110001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001100110001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011001100110010000) && ({row_reg, col_reg}<19'b0011001101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001101001010001) && ({row_reg, col_reg}<19'b0011001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011001101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011001101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011001110000000000) && ({row_reg, col_reg}<19'b0011001110010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001110010010101) && ({row_reg, col_reg}<19'b0011001110010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110010010111) && ({row_reg, col_reg}<19'b0011001110010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001110010110011) && ({row_reg, col_reg}<19'b0011001110010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001110010110110) && ({row_reg, col_reg}<19'b0011001110010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110010111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001110010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110010111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001110010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110010111111) && ({row_reg, col_reg}<19'b0011001110011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110011010001) && ({row_reg, col_reg}<19'b0011001110011010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110011010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110011010100) && ({row_reg, col_reg}<19'b0011001110011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110011010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001110011010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011001110011011000) && ({row_reg, col_reg}<19'b0011001110011100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110011100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011001110011100010) && ({row_reg, col_reg}<19'b0011001110011100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110011100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001110011100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011001110011100110) && ({row_reg, col_reg}<19'b0011001110011101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110011101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001110011101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001110011101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001110011101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001110011101100) && ({row_reg, col_reg}<19'b0011001110011101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110011101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011001110011101111) && ({row_reg, col_reg}<19'b0011001110011110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001110011110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001110011110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011001110011110011) && ({row_reg, col_reg}<19'b0011001110011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110011110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001110011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110011111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110011111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001110011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110011111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001110011111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110011111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011001110100000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110100000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001110100000010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011001110100000011) && ({row_reg, col_reg}<19'b0011001110100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001110100000101) && ({row_reg, col_reg}<19'b0011001110100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110100000111) && ({row_reg, col_reg}<19'b0011001110100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110100010001) && ({row_reg, col_reg}<19'b0011001110100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110100010100) && ({row_reg, col_reg}<19'b0011001110100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110100010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011001110100010111) && ({row_reg, col_reg}<19'b0011001110100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110100011010) && ({row_reg, col_reg}<19'b0011001110100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001110100011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001110100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110100100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011001110100100010) && ({row_reg, col_reg}<19'b0011001110100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001110100101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001110100101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001110100101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001110100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110100101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001110100101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001110100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001110100110001) && ({row_reg, col_reg}<19'b0011001110100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110100110011) && ({row_reg, col_reg}<19'b0011001110100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110100111001) && ({row_reg, col_reg}<19'b0011001110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001110100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011001110100111111) && ({row_reg, col_reg}<19'b0011001110101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001110101000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011001110101000011) && ({row_reg, col_reg}<19'b0011001110101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110101000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011001110101000110) && ({row_reg, col_reg}<19'b0011001110101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011001110101001000) && ({row_reg, col_reg}<19'b0011001110101001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001110101001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001110101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110101001100) && ({row_reg, col_reg}<19'b0011001110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001110101001111) && ({row_reg, col_reg}<19'b0011001110101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011001110101010001) && ({row_reg, col_reg}<19'b0011001110101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001110101010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001110101010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110101011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001110101011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011001110101011010) && ({row_reg, col_reg}<19'b0011001110101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110101011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001110101011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001110101011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001110101011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011001110101100000) && ({row_reg, col_reg}<19'b0011001110101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001110101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110101100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001110101100100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001110101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110101100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001110101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001110101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001110101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011001110101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110101101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001110101101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011001110101101111) && ({row_reg, col_reg}<19'b0011001110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110101111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001110101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001110101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110101111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011001110101111100) && ({row_reg, col_reg}<19'b0011001110101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110101111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011001110101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001110110000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011001110110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001110110000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011001110110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110110000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001110110000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001110110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001110110001000) && ({row_reg, col_reg}<19'b0011001110110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110110001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001110110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011001110110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011001110110001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011001110110001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011001110110001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011001110110010000) && ({row_reg, col_reg}<19'b0011001111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011001111001010001) && ({row_reg, col_reg}<19'b0011001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011001111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011001111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011010000000000000) && ({row_reg, col_reg}<19'b0011010000010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010000010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010000010110011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000010110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011010000010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010000010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010000010111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010000010111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010000010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010000010111110) && ({row_reg, col_reg}<19'b0011010000011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011010000011011000) && ({row_reg, col_reg}<19'b0011010000011011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010000011011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010000011011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010000011011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011010000011011111) && ({row_reg, col_reg}<19'b0011010000011100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010000011100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011010000011100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010000011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000011100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000011100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010000011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000011100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010000011101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010000011101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000011101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000011101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010000011101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010000011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010000011101110) && ({row_reg, col_reg}<19'b0011010000011110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010000011110000) && ({row_reg, col_reg}<19'b0011010000011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000011111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010000011111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010000011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000011111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011010000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010000100000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010000100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010000100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010000100000100) && ({row_reg, col_reg}<19'b0011010000100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010000100010001) && ({row_reg, col_reg}<19'b0011010000100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010000100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010000100010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010000100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000100011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010000100011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010000100011010) && ({row_reg, col_reg}<19'b0011010000100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011010000100011100) && ({row_reg, col_reg}<19'b0011010000100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010000100011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010000100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000100100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011010000100100001) && ({row_reg, col_reg}<19'b0011010000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010000100100110) && ({row_reg, col_reg}<19'b0011010000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010000100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000100101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010000100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010000100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010000100101110) && ({row_reg, col_reg}<19'b0011010000100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000100110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011010000100110001) && ({row_reg, col_reg}<19'b0011010000100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010000100110100) && ({row_reg, col_reg}<19'b0011010000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010000100110111) && ({row_reg, col_reg}<19'b0011010000100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010000100111010) && ({row_reg, col_reg}<19'b0011010000100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010000100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010000100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010000101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010000101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010000101000101) && ({row_reg, col_reg}<19'b0011010000101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010000101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010000101010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010000101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000101010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011010000101010110) && ({row_reg, col_reg}<19'b0011010000101011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010000101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010000101011010) && ({row_reg, col_reg}<19'b0011010000101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000101011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000101011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000101011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000101011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011010000101100000) && ({row_reg, col_reg}<19'b0011010000101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000101100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010000101100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000101100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011010000101101000) && ({row_reg, col_reg}<19'b0011010000101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000101101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010000101101101) && ({row_reg, col_reg}<19'b0011010000101101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000101101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010000101110000) && ({row_reg, col_reg}<19'b0011010000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000101111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010000101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010000101111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010000101111100) && ({row_reg, col_reg}<19'b0011010000101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000101111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010000110000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011010000110000001) && ({row_reg, col_reg}<19'b0011010000110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000110000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011010000110000100) && ({row_reg, col_reg}<19'b0011010000110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000110001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011010000110001001) && ({row_reg, col_reg}<19'b0011010000110001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000110001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010000110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010000110001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000110001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010000110001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010000110010000) && ({row_reg, col_reg}<19'b0011010001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011010001001010001) && ({row_reg, col_reg}<19'b0011010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011010001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011010001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011010010000000000) && ({row_reg, col_reg}<19'b0011010010010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010010010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010010110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010010010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010010110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010010010110111) && ({row_reg, col_reg}<19'b0011010010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010010111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010010111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010010010111100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010010010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010010010111110) && ({row_reg, col_reg}<19'b0011010010011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011010010011011000) && ({row_reg, col_reg}<19'b0011010010011011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010010011011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010010011011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010010011011110) && ({row_reg, col_reg}<19'b0011010010011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010011100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010010011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010011100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011010010011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010011100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010010011100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010010011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010011100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010010011101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011010010011101001) && ({row_reg, col_reg}<19'b0011010010011101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010010011101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011010010011101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010010011101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010010011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010010011110000) && ({row_reg, col_reg}<19'b0011010010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010011111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010010011111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010010011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010011111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011010010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010100000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010010100000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010010100000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010010100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010010100000100) && ({row_reg, col_reg}<19'b0011010010100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010010100000111) && ({row_reg, col_reg}<19'b0011010010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010010100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011010010100010010) && ({row_reg, col_reg}<19'b0011010010100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010010100010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010010100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010100011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011010010100011001) && ({row_reg, col_reg}<19'b0011010010100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010100011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010100100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011010010100100001) && ({row_reg, col_reg}<19'b0011010010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010010100100110) && ({row_reg, col_reg}<19'b0011010010100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010010100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010100101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010010100101110) && ({row_reg, col_reg}<19'b0011010010100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010100110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011010010100110001) && ({row_reg, col_reg}<19'b0011010010100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010010100110100) && ({row_reg, col_reg}<19'b0011010010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010010100110111) && ({row_reg, col_reg}<19'b0011010010100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010010100111010) && ({row_reg, col_reg}<19'b0011010010100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010010100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010010101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010010101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010010101000101) && ({row_reg, col_reg}<19'b0011010010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010010101010001) && ({row_reg, col_reg}<19'b0011010010101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010101010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010101010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010101010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010101010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011010010101011000) && ({row_reg, col_reg}<19'b0011010010101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010101011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010010101011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010010101011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010101011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010010101011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010010101100000) && ({row_reg, col_reg}<19'b0011010010101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010010101100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010010101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010101100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011010010101101000) && ({row_reg, col_reg}<19'b0011010010101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010101101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010010101101101) && ({row_reg, col_reg}<19'b0011010010101101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010101101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010010101110000) && ({row_reg, col_reg}<19'b0011010010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010101111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010010101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010101111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010010101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010010101111100) && ({row_reg, col_reg}<19'b0011010010101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010010101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010110000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010010110000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010010110000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010010110000100) && ({row_reg, col_reg}<19'b0011010010110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010110001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010010110001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010010110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010110001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010010110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010010110001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010110001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010010110001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011010010110010000) && ({row_reg, col_reg}<19'b0011010011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011010011001010001) && ({row_reg, col_reg}<19'b0011010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011010011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011010011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011010100000000000) && ({row_reg, col_reg}<19'b0011010100010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010100010110001) && ({row_reg, col_reg}<19'b0011010100010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100010110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010100010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100010110101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010100010110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010100010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100010111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011010100010111011) && ({row_reg, col_reg}<19'b0011010100010111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010100010111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010100010111110) && ({row_reg, col_reg}<19'b0011010100011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100011100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010100011100011) && ({row_reg, col_reg}<19'b0011010100011100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010100011100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010100011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100011100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010100011101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010100011101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010100011101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010100011101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010100011101100) && ({row_reg, col_reg}<19'b0011010100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100011111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010100011111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010100011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100011111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010100100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100100000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010100100000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010100100000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010100100000100) && ({row_reg, col_reg}<19'b0011010100100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010100100000111) && ({row_reg, col_reg}<19'b0011010100100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010100100010011) && ({row_reg, col_reg}<19'b0011010100100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100100010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100100010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010100100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010100100011001) && ({row_reg, col_reg}<19'b0011010100100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010100100011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100100100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010100100100001) && ({row_reg, col_reg}<19'b0011010100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010100100100110) && ({row_reg, col_reg}<19'b0011010100100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010100100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100100101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010100100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010100100101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010100100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100100110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011010100100110001) && ({row_reg, col_reg}<19'b0011010100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010100100110100) && ({row_reg, col_reg}<19'b0011010100100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010100100110111) && ({row_reg, col_reg}<19'b0011010100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010100100111010) && ({row_reg, col_reg}<19'b0011010100100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010100100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010100100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010100101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010100101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010100101000101) && ({row_reg, col_reg}<19'b0011010100101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100101010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010100101010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010100101010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100101010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011010100101011000) && ({row_reg, col_reg}<19'b0011010100101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100101011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010100101011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010100101011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100101011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010100101011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011010100101011111) && ({row_reg, col_reg}<19'b0011010100101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010100101100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010100101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100101100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011010100101101000) && ({row_reg, col_reg}<19'b0011010100101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100101101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010100101101101) && ({row_reg, col_reg}<19'b0011010100101101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100101101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010100101110000) && ({row_reg, col_reg}<19'b0011010100101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100101111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010100101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100101111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010100101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010100101111100) && ({row_reg, col_reg}<19'b0011010100101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100101111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010100101111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010100110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010100110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010100110000011) && ({row_reg, col_reg}<19'b0011010100110001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010100110001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010100110001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010100110001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011010100110001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010100110001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010100110001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010100110001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011010100110010000) && ({row_reg, col_reg}<19'b0011010101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011010101001010001) && ({row_reg, col_reg}<19'b0011010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011010101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011010101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011010110000000000) && ({row_reg, col_reg}<19'b0011010110010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110010110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010110010110001) && ({row_reg, col_reg}<19'b0011010110010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110010110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110010110101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010110010110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011010110010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110010111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011010110010111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010110010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110010111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011010110010111110) && ({row_reg, col_reg}<19'b0011010110011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110011100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110011100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010110011100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010110011100110) && ({row_reg, col_reg}<19'b0011010110011101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010110011101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010110011101011) && ({row_reg, col_reg}<19'b0011010110011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110011101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010110011110000) && ({row_reg, col_reg}<19'b0011010110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110011111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010110011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110011111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110100000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010110100000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010110100000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110100000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010110100000100) && ({row_reg, col_reg}<19'b0011010110100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010110100000111) && ({row_reg, col_reg}<19'b0011010110100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011010110100010001) && ({row_reg, col_reg}<19'b0011010110100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010110100010011) && ({row_reg, col_reg}<19'b0011010110100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010110100010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110100010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010110100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010110100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110100011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110100011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010110100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011010110100100001) && ({row_reg, col_reg}<19'b0011010110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010110100100110) && ({row_reg, col_reg}<19'b0011010110100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010110100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110100101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011010110100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011010110100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110100101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010110100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110100110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010110100110100) && ({row_reg, col_reg}<19'b0011010110100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010110100110111) && ({row_reg, col_reg}<19'b0011010110100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010110100111010) && ({row_reg, col_reg}<19'b0011010110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010110100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010110100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010110101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010110101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011010110101000101) && ({row_reg, col_reg}<19'b0011010110101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110101010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010110101010111) && ({row_reg, col_reg}<19'b0011010110101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110101011010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011010110101011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011010110101011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110101011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010110101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010110101011111) && ({row_reg, col_reg}<19'b0011010110101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011010110101100011) && ({row_reg, col_reg}<19'b0011010110101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110101100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010110101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110101100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011010110101101000) && ({row_reg, col_reg}<19'b0011010110101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110101101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010110101101101) && ({row_reg, col_reg}<19'b0011010110101101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110101101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011010110101110000) && ({row_reg, col_reg}<19'b0011010110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110101111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010110101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110101111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010110101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010110101111100) && ({row_reg, col_reg}<19'b0011010110101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110101111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011010110101111111) && ({row_reg, col_reg}<19'b0011010110110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110110000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011010110110000010) && ({row_reg, col_reg}<19'b0011010110110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110110000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011010110110000101) && ({row_reg, col_reg}<19'b0011010110110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110110000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011010110110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011010110110001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010110110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110110001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010110110001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010110110001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011010110110001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010110110001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010110110010000) && ({row_reg, col_reg}<19'b0011010111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011010111001010001) && ({row_reg, col_reg}<19'b0011010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011010111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011010111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011011000000000000) && ({row_reg, col_reg}<19'b0011011000010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011000010110001) && ({row_reg, col_reg}<19'b0011011000010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000010110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011000010110100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011000010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000010110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011000010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000010111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011000010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000010111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011000010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011000010111111) && ({row_reg, col_reg}<19'b0011011000011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000011100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011000011100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011000011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000011100100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011000011100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011000011100110) && ({row_reg, col_reg}<19'b0011011000011101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011000011101000) && ({row_reg, col_reg}<19'b0011011000011101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000011101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011000011101100) && ({row_reg, col_reg}<19'b0011011000011101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011000011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000011101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011000011110000) && ({row_reg, col_reg}<19'b0011011000011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000011111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011000011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000011111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011000011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011000011111111) && ({row_reg, col_reg}<19'b0011011000100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011000100000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000100000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011011000100000100) && ({row_reg, col_reg}<19'b0011011000100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011000100000111) && ({row_reg, col_reg}<19'b0011011000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011000100010001) && ({row_reg, col_reg}<19'b0011011000100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000100010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011000100010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000100010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011011000100011000) && ({row_reg, col_reg}<19'b0011011000100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000100011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000100011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011000100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011000100100011) && ({row_reg, col_reg}<19'b0011011000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011000100100110) && ({row_reg, col_reg}<19'b0011011000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011000100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000100101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011011000100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011000100101100) && ({row_reg, col_reg}<19'b0011011000100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100101110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011000100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000100110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011000100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011000100110100) && ({row_reg, col_reg}<19'b0011011000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011000100110111) && ({row_reg, col_reg}<19'b0011011000100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011000100111010) && ({row_reg, col_reg}<19'b0011011000100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011000100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011000100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011000101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011000101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011000101000101) && ({row_reg, col_reg}<19'b0011011000101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011000101010010) && ({row_reg, col_reg}<19'b0011011000101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011000101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000101010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011000101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011011000101011011) && ({row_reg, col_reg}<19'b0011011000101011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000101011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011011000101011110) && ({row_reg, col_reg}<19'b0011011000101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011000101100011) && ({row_reg, col_reg}<19'b0011011000101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011000101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000101100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011011000101101000) && ({row_reg, col_reg}<19'b0011011000101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011000101101101) && ({row_reg, col_reg}<19'b0011011000101101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000101101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011000101110000) && ({row_reg, col_reg}<19'b0011011000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011000101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011000101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011000101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000110000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011000110000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011000110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000110000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011000110000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011000110000101) && ({row_reg, col_reg}<19'b0011011000110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011000110000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011000110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011000110001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011011000110001010) && ({row_reg, col_reg}<19'b0011011000110001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000110001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011000110001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011000110001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011011000110010000) && ({row_reg, col_reg}<19'b0011011001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011001001010001) && ({row_reg, col_reg}<19'b0011011001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011011001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011011001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011011010000000000) && ({row_reg, col_reg}<19'b0011011010010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011010010110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011010010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010010110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011010010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011010010111000) && ({row_reg, col_reg}<19'b0011011010010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010010111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011011010010111100) && ({row_reg, col_reg}<19'b0011011010010111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011010010111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011011010010111111) && ({row_reg, col_reg}<19'b0011011010011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011010011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010011100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011011010011100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011010011100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011010011100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011010011100101) && ({row_reg, col_reg}<19'b0011011010011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010011100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010011101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011010011101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011010011101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010011101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011010011101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011010011101110) && ({row_reg, col_reg}<19'b0011011010011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010011111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011011010011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010011111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011010011111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011010011111111) && ({row_reg, col_reg}<19'b0011011010100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011010100000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011010100000100) && ({row_reg, col_reg}<19'b0011011010100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011010100000111) && ({row_reg, col_reg}<19'b0011011010100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011011010100010101) && ({row_reg, col_reg}<19'b0011011010100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010100010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011010100011000) && ({row_reg, col_reg}<19'b0011011010100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011010100011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011010100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011010100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011011010100100001) && ({row_reg, col_reg}<19'b0011011010100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011010100100011) && ({row_reg, col_reg}<19'b0011011010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011010100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011010100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011010100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010100101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011010100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011010100101100) && ({row_reg, col_reg}<19'b0011011010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100101110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011010100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010100110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011010100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011010100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011010100110100) && ({row_reg, col_reg}<19'b0011011010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011010100110111) && ({row_reg, col_reg}<19'b0011011010100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011010100111010) && ({row_reg, col_reg}<19'b0011011010100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011010100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011010100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011010101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011010101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011010101000101) && ({row_reg, col_reg}<19'b0011011010101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011010101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011011010101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011010101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010101010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011010101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011010101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011010101011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011010101011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011010101011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011010101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011010101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011010101100000) && ({row_reg, col_reg}<19'b0011011010101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011010101100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011010101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010101100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011011010101101000) && ({row_reg, col_reg}<19'b0011011010101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011010101101101) && ({row_reg, col_reg}<19'b0011011010101101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010101101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011010101110000) && ({row_reg, col_reg}<19'b0011011010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011010101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010101111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011011010101111011) && ({row_reg, col_reg}<19'b0011011010101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010101111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011010101111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011010101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011010110000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011010110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011010110000011) && ({row_reg, col_reg}<19'b0011011010110000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011010110000101) && ({row_reg, col_reg}<19'b0011011010110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010110000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011010110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011010110001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011010110001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011010110001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011010110001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011010110001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011010110001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011010110001111) && ({row_reg, col_reg}<19'b0011011011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011011001010001) && ({row_reg, col_reg}<19'b0011011011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011011011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011011011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011011100000000000) && ({row_reg, col_reg}<19'b0011011100010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011100010110010) && ({row_reg, col_reg}<19'b0011011100010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100010110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011100010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100010110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011100010110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011100010111000) && ({row_reg, col_reg}<19'b0011011100010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100010111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011100010111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100010111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011011100010111111) && ({row_reg, col_reg}<19'b0011011100011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011100011011010) && ({row_reg, col_reg}<19'b0011011100011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011100011011110) && ({row_reg, col_reg}<19'b0011011100011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100011100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011100011100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011100011100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011100011100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011011100011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100011100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100011101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011100011101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100011101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100011101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100011101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011100011101110) && ({row_reg, col_reg}<19'b0011011100011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100011111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011100011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100011111101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011100011111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011100011111111) && ({row_reg, col_reg}<19'b0011011100100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011100100000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100100000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011100100000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011100100000101) && ({row_reg, col_reg}<19'b0011011100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011100100010001) && ({row_reg, col_reg}<19'b0011011100100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011011100100010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011100100010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100100010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011011100100010111) && ({row_reg, col_reg}<19'b0011011100100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100100011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011100100011011) && ({row_reg, col_reg}<19'b0011011100100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100100011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011100100011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011100100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011011100100100001) && ({row_reg, col_reg}<19'b0011011100100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011100100100011) && ({row_reg, col_reg}<19'b0011011100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011100100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100100101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011100100101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011100100101100) && ({row_reg, col_reg}<19'b0011011100100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011100100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100100110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011100100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011100100110111) && ({row_reg, col_reg}<19'b0011011100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011100100111010) && ({row_reg, col_reg}<19'b0011011100100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011100100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011100100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011100101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011100101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011100101000101) && ({row_reg, col_reg}<19'b0011011100101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100101010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011100101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100101010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011100101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011100101010111) && ({row_reg, col_reg}<19'b0011011100101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100101011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011100101011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011100101011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011100101011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011100101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011100101100000) && ({row_reg, col_reg}<19'b0011011100101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100101100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011100101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100101100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011011100101101000) && ({row_reg, col_reg}<19'b0011011100101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100101101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011100101101101) && ({row_reg, col_reg}<19'b0011011100101101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100101101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011100101110000) && ({row_reg, col_reg}<19'b0011011100101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100101111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011100101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011011100101111011) && ({row_reg, col_reg}<19'b0011011100101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100101111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011100101111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011100101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100110000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011011100110000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011100110000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011100110000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011100110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011100110000110) && ({row_reg, col_reg}<19'b0011011100110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011100110001010) && ({row_reg, col_reg}<19'b0011011100110001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011100110001100) && ({row_reg, col_reg}<19'b0011011101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011101001010001) && ({row_reg, col_reg}<19'b0011011101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011011101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011011101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011011110000000000) && ({row_reg, col_reg}<19'b0011011110010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011110010110010) && ({row_reg, col_reg}<19'b0011011110010110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110010110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011011110010110101) && ({row_reg, col_reg}<19'b0011011110010110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110010110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011110010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011110010111010) && ({row_reg, col_reg}<19'b0011011110010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110010111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011110010111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110010111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011011110010111111) && ({row_reg, col_reg}<19'b0011011110011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011110011011000) && ({row_reg, col_reg}<19'b0011011110011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011110011011010) && ({row_reg, col_reg}<19'b0011011110011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110011100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011110011100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011011110011100010) && ({row_reg, col_reg}<19'b0011011110011100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110011100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011110011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110011100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011110011100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110011101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011011110011101010) && ({row_reg, col_reg}<19'b0011011110011101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110011101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011110011101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011011110011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110011101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011110011110000) && ({row_reg, col_reg}<19'b0011011110011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110011111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011110011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110011111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011110011111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011110011111111) && ({row_reg, col_reg}<19'b0011011110100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011110100000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011110100000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011110100000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011110100000101) && ({row_reg, col_reg}<19'b0011011110100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011110100010001) && ({row_reg, col_reg}<19'b0011011110100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011110100010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011110100010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110100010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011110100010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110100011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011110100011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011110100011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011011110100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110100011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110100011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011110100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011011110100100001) && ({row_reg, col_reg}<19'b0011011110100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011110100100011) && ({row_reg, col_reg}<19'b0011011110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110100101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011110100101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011110100101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011011110100101100) && ({row_reg, col_reg}<19'b0011011110100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011110100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110100110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011110100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011110100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011110100110111) && ({row_reg, col_reg}<19'b0011011110100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011110100111010) && ({row_reg, col_reg}<19'b0011011110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011110100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011110100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011011110101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011110101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011110101000101) && ({row_reg, col_reg}<19'b0011011110101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110101010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110101010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011110101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011011110101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110101011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011110101011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011110101011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011011110101011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011110101011110) && ({row_reg, col_reg}<19'b0011011110101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110101100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011011110101100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011011110101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110101100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011011110101101000) && ({row_reg, col_reg}<19'b0011011110101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110101101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011011110101101101) && ({row_reg, col_reg}<19'b0011011110101101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110101101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011110101110000) && ({row_reg, col_reg}<19'b0011011110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011110101111000) && ({row_reg, col_reg}<19'b0011011110101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110101111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011011110101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110101111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011011110101111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011110101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110110000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011011110110000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011110110000010) && ({row_reg, col_reg}<19'b0011011110110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110110000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011110110000110) && ({row_reg, col_reg}<19'b0011011110110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110110001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011011110110001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011011110110001010) && ({row_reg, col_reg}<19'b0011011110110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011011110110001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011011110110001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011011110110010000) && ({row_reg, col_reg}<19'b0011011111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011011111001010001) && ({row_reg, col_reg}<19'b0011011111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011011111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011011111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011100000000000000) && ({row_reg, col_reg}<19'b0011100000010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100000010110001) && ({row_reg, col_reg}<19'b0011100000010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100000010110011) && ({row_reg, col_reg}<19'b0011100000010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000010110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100000010110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000010110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100000010111000) && ({row_reg, col_reg}<19'b0011100000010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100000010111010) && ({row_reg, col_reg}<19'b0011100000010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000010111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011100000010111101) && ({row_reg, col_reg}<19'b0011100000010111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100000010111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011100000011000000) && ({row_reg, col_reg}<19'b0011100000011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100000011000111) && ({row_reg, col_reg}<19'b0011100000011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100000011001001) && ({row_reg, col_reg}<19'b0011100000011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100000011001110) && ({row_reg, col_reg}<19'b0011100000011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100000011010010) && ({row_reg, col_reg}<19'b0011100000011010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000011010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100000011011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100000011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100000011011010) && ({row_reg, col_reg}<19'b0011100000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100000011011101) && ({row_reg, col_reg}<19'b0011100000011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100000011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000011100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100000011100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100000011100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000011100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011100000011100100) && ({row_reg, col_reg}<19'b0011100000011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000011100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100000011100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000011101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011100000011101010) && ({row_reg, col_reg}<19'b0011100000011101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000011101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100000011101101) && ({row_reg, col_reg}<19'b0011100000011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100000011110000) && ({row_reg, col_reg}<19'b0011100000011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000011111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011100000011111001) && ({row_reg, col_reg}<19'b0011100000011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000011111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100000011111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100000011111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000011111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011100000011111111) && ({row_reg, col_reg}<19'b0011100000100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000100000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011100000100000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000100000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100000100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100000100000101) && ({row_reg, col_reg}<19'b0011100000100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000100010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000100010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000100010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100000100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100000100010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100000100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000100011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100000100011011) && ({row_reg, col_reg}<19'b0011100000100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000100011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011100000100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100000100100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100000100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100000100100100) && ({row_reg, col_reg}<19'b0011100000100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100000100100110) && ({row_reg, col_reg}<19'b0011100000100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100000100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100000100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100000100101011) && ({row_reg, col_reg}<19'b0011100000100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100000100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100000100110001) && ({row_reg, col_reg}<19'b0011100000100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100000100110110) && ({row_reg, col_reg}<19'b0011100000100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100000100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011100000100111111) && ({row_reg, col_reg}<19'b0011100000101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100000101000010) && ({row_reg, col_reg}<19'b0011100000101000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100000101000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100000101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100000101000111) && ({row_reg, col_reg}<19'b0011100000101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100000101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000101010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100000101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100000101010111) && ({row_reg, col_reg}<19'b0011100000101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000101011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100000101011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100000101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100000101011111) && ({row_reg, col_reg}<19'b0011100000101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100000101100010) && ({row_reg, col_reg}<19'b0011100000101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100000101100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100000101100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100000101100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100000101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011100000101101010) && ({row_reg, col_reg}<19'b0011100000101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100000101101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000101101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100000101101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100000101110000) && ({row_reg, col_reg}<19'b0011100000101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100000101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100000101111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100000101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000101111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011100000101111011) && ({row_reg, col_reg}<19'b0011100000101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100000101111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000101111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100000110000000) && ({row_reg, col_reg}<19'b0011100000110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100000110110000) && ({row_reg, col_reg}<19'b0011100000110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011100000110110011) && ({row_reg, col_reg}<19'b0011100000110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100000110111000) && ({row_reg, col_reg}<19'b0011100000110111011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0011100000110111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100000110111100) && ({row_reg, col_reg}<19'b0011100000111000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011100000111000000) && ({row_reg, col_reg}<19'b0011100001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100001001010001) && ({row_reg, col_reg}<19'b0011100001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011100001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011100001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011100010000000000) && ({row_reg, col_reg}<19'b0011100010010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100010010110001) && ({row_reg, col_reg}<19'b0011100010010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010010110011) && ({row_reg, col_reg}<19'b0011100010010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010010110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100010010110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100010010110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100010010111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100010010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100010010111010) && ({row_reg, col_reg}<19'b0011100010010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010010111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100010010111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100010010111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100010010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010011000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100010011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010011000010) && ({row_reg, col_reg}<19'b0011100010011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010011000110) && ({row_reg, col_reg}<19'b0011100010011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100010011001110) && ({row_reg, col_reg}<19'b0011100010011010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010011010010) && ({row_reg, col_reg}<19'b0011100010011011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100010011011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100010011011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100010011011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100010011011110) && ({row_reg, col_reg}<19'b0011100010011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010011100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100010011100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100010011100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100010011100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011100010011100100) && ({row_reg, col_reg}<19'b0011100010011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010011100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010011100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010011101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011100010011101010) && ({row_reg, col_reg}<19'b0011100010011101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010011101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010011101101) && ({row_reg, col_reg}<19'b0011100010011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010011110000) && ({row_reg, col_reg}<19'b0011100010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100010011111001) && ({row_reg, col_reg}<19'b0011100010011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010011111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100010011111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100010011111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010011111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100010011111111) && ({row_reg, col_reg}<19'b0011100010100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010100000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011100010100000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010100000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100010100000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100010100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100010100000110) && ({row_reg, col_reg}<19'b0011100010100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010100001000) && ({row_reg, col_reg}<19'b0011100010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010100010001) && ({row_reg, col_reg}<19'b0011100010100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010100010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100010100010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010100010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100010100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100010100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010100011000) && ({row_reg, col_reg}<19'b0011100010100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010100011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100010100011011) && ({row_reg, col_reg}<19'b0011100010100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010100011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100010100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100010100100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100010100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100010100100100) && ({row_reg, col_reg}<19'b0011100010100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100010100100110) && ({row_reg, col_reg}<19'b0011100010100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100010100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100010100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100010100101011) && ({row_reg, col_reg}<19'b0011100010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100010100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100010100110001) && ({row_reg, col_reg}<19'b0011100010100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100010100110110) && ({row_reg, col_reg}<19'b0011100010100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100010100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011100010100111111) && ({row_reg, col_reg}<19'b0011100010101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100010101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100010101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010101000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100010101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010101000111) && ({row_reg, col_reg}<19'b0011100010101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100010101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010101010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100010101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100010101010111) && ({row_reg, col_reg}<19'b0011100010101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010101011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100010101011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100010101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010101011111) && ({row_reg, col_reg}<19'b0011100010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100010101100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100010101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010101100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011100010101100111) && ({row_reg, col_reg}<19'b0011100010101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011100010101101010) && ({row_reg, col_reg}<19'b0011100010101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100010101101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010101101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100010101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100010101110000) && ({row_reg, col_reg}<19'b0011100010101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100010101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100010101111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100010101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010101111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100010101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100010101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100010101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010101111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011100010110000000) && ({row_reg, col_reg}<19'b0011100010110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100010110110000) && ({row_reg, col_reg}<19'b0011100010110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011100010110110011) && ({row_reg, col_reg}<19'b0011100010110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100010110110111) && ({row_reg, col_reg}<19'b0011100010110111010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0011100010110111010) && ({row_reg, col_reg}<19'b0011100010110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100010110111100) && ({row_reg, col_reg}<19'b0011100010110111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011100010110111110) && ({row_reg, col_reg}<19'b0011100010111000000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0011100010111000000) && ({row_reg, col_reg}<19'b0011100011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100011001010001) && ({row_reg, col_reg}<19'b0011100011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011100011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011100011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011100100000000000) && ({row_reg, col_reg}<19'b0011100100010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100010110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100100010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100100010110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100010111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100100010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100100010111010) && ({row_reg, col_reg}<19'b0011100100010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100010111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100100010111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100100010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100011000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100100011000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011100100011000010) && ({row_reg, col_reg}<19'b0011100100011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100100011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100100011000111) && ({row_reg, col_reg}<19'b0011100100011011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100100011011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100100011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100100011011101) && ({row_reg, col_reg}<19'b0011100100011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100100011100000) && ({row_reg, col_reg}<19'b0011100100011100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100100011100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100100011100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100100011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100011100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100100011100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100100011100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100011101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100100011101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100100011101010) && ({row_reg, col_reg}<19'b0011100100011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100100011110000) && ({row_reg, col_reg}<19'b0011100100011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100011111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011100100011111101) && ({row_reg, col_reg}<19'b0011100100011111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011100100100000010) && ({row_reg, col_reg}<19'b0011100100100000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100100000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100100100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100100100000110) && ({row_reg, col_reg}<19'b0011100100100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100100100001000) && ({row_reg, col_reg}<19'b0011100100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100100100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100100100010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100100100010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100100010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100100100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100100100010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011100100100011000) && ({row_reg, col_reg}<19'b0011100100100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100100011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011100100100011011) && ({row_reg, col_reg}<19'b0011100100100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100100100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100100100100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100100100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100100100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100100100100100) && ({row_reg, col_reg}<19'b0011100100100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100100100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100100100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100100100101011) && ({row_reg, col_reg}<19'b0011100100100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100100100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100100100110001) && ({row_reg, col_reg}<19'b0011100100100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100100100110110) && ({row_reg, col_reg}<19'b0011100100100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100100100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011100100100111111) && ({row_reg, col_reg}<19'b0011100100101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100100101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100100101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100101000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011100100101000101) && ({row_reg, col_reg}<19'b0011100100101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100100101010011) && ({row_reg, col_reg}<19'b0011100100101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100100101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100100101010111) && ({row_reg, col_reg}<19'b0011100100101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100100101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100101011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100100101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100100101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100100101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100100101100001) && ({row_reg, col_reg}<19'b0011100100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100100101100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100100101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100101100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011100100101100111) && ({row_reg, col_reg}<19'b0011100100101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011100100101101010) && ({row_reg, col_reg}<19'b0011100100101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100100101101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100101101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100100101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100100101110000) && ({row_reg, col_reg}<19'b0011100100101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100100101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100100101111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100100101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100101111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100100101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100100101111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100100101111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100101111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011100100110000000) && ({row_reg, col_reg}<19'b0011100100110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100100110110000) && ({row_reg, col_reg}<19'b0011100100110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011100100110110011) && ({row_reg, col_reg}<19'b0011100100110110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100100110110111) && ({row_reg, col_reg}<19'b0011100100110111010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0011100100110111010) && ({row_reg, col_reg}<19'b0011100100110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100100110111101) && ({row_reg, col_reg}<19'b0011100100110111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0011100100110111111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0011100100111000000) && ({row_reg, col_reg}<19'b0011100101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100101001010001) && ({row_reg, col_reg}<19'b0011100101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011100101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011100101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011100110000000000) && ({row_reg, col_reg}<19'b0011100110010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100110010110001) && ({row_reg, col_reg}<19'b0011100110010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100110010110100) && ({row_reg, col_reg}<19'b0011100110010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110010110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011100110010110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110010111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100110010111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011100110010111010) && ({row_reg, col_reg}<19'b0011100110010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011100110010111111) && ({row_reg, col_reg}<19'b0011100110011000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110011000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100110011000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011100110011000011) && ({row_reg, col_reg}<19'b0011100110011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110011000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100110011000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100110011001000) && ({row_reg, col_reg}<19'b0011100110011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100110011001101) && ({row_reg, col_reg}<19'b0011100110011010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100110011010011) && ({row_reg, col_reg}<19'b0011100110011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100110011011000) && ({row_reg, col_reg}<19'b0011100110011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110011011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100110011011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100110011100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110011100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100110011100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011100110011100011) && ({row_reg, col_reg}<19'b0011100110011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110011100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011100110011100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100110011100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110011101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110011101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100110011101010) && ({row_reg, col_reg}<19'b0011100110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100110011111001) && ({row_reg, col_reg}<19'b0011100110011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100110011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100110011111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100110011111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110011111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100110100000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100110100000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011100110100000101) && ({row_reg, col_reg}<19'b0011100110100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011100110100001000) && ({row_reg, col_reg}<19'b0011100110100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100110100010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011100110100010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100110100010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110100010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100110100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011100110100011000) && ({row_reg, col_reg}<19'b0011100110100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110100011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011100110100011011) && ({row_reg, col_reg}<19'b0011100110100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100110100011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100110100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100110100100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100110100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100110100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100110100100100) && ({row_reg, col_reg}<19'b0011100110100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100110100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100110100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100110100101011) && ({row_reg, col_reg}<19'b0011100110100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100110100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100110100110001) && ({row_reg, col_reg}<19'b0011100110100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011100110100110110) && ({row_reg, col_reg}<19'b0011100110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100110100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011100110100111111) && ({row_reg, col_reg}<19'b0011100110101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100110101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011100110101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100110101000101) && ({row_reg, col_reg}<19'b0011100110101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100110101010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011100110101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011100110101010101) && ({row_reg, col_reg}<19'b0011100110101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100110101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110101011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011100110101011100) && ({row_reg, col_reg}<19'b0011100110101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100110101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011100110101100001) && ({row_reg, col_reg}<19'b0011100110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110101100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110101100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100110101100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011100110101100111) && ({row_reg, col_reg}<19'b0011100110101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011100110101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100110101101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100110101101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110101101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011100110101101111) && ({row_reg, col_reg}<19'b0011100110101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011100110101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011100110101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011100110101111010) && ({row_reg, col_reg}<19'b0011100110101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110101111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011100110101111101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110101111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011100110110000000) && ({row_reg, col_reg}<19'b0011100110110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100110110110000) && ({row_reg, col_reg}<19'b0011100110110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011100110110110011) && ({row_reg, col_reg}<19'b0011100110110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011100110110111000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0011100110110111001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0011100110110111010) && ({row_reg, col_reg}<19'b0011100110110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100110110111110) && ({row_reg, col_reg}<19'b0011100110111000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011100110111000000) && ({row_reg, col_reg}<19'b0011100111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011100111001010001) && ({row_reg, col_reg}<19'b0011100111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011100111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011100111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011101000000000000) && ({row_reg, col_reg}<19'b0011101000010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101000010110001) && ({row_reg, col_reg}<19'b0011101000010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101000010110100) && ({row_reg, col_reg}<19'b0011101000010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000010110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101000010110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101000010111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000010111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101000010111010) && ({row_reg, col_reg}<19'b0011101000010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101000010111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011101000011000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000011000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101000011000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101000011000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101000011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101000011000101) && ({row_reg, col_reg}<19'b0011101000011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101000011001000) && ({row_reg, col_reg}<19'b0011101000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000011011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101000011011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101000011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000011100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101000011100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101000011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101000011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101000011100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101000011100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101000011100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000011101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011101000011101001) && ({row_reg, col_reg}<19'b0011101000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101000011111001) && ({row_reg, col_reg}<19'b0011101000011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101000011111011) && ({row_reg, col_reg}<19'b0011101000011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000011111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101000011111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000011111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011101000100000000) && ({row_reg, col_reg}<19'b0011101000100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101000100000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101000100000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000100000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011101000100000101) && ({row_reg, col_reg}<19'b0011101000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000100010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101000100010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101000100010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000100010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011101000100010101) && ({row_reg, col_reg}<19'b0011101000100010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000100010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101000100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000100011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101000100011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011101000100011011) && ({row_reg, col_reg}<19'b0011101000100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101000100011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011101000100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101000100100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101000100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101000100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101000100100100) && ({row_reg, col_reg}<19'b0011101000100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101000100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101000100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101000100101011) && ({row_reg, col_reg}<19'b0011101000100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101000100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101000100110001) && ({row_reg, col_reg}<19'b0011101000100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101000100110110) && ({row_reg, col_reg}<19'b0011101000100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101000100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011101000100111111) && ({row_reg, col_reg}<19'b0011101000101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101000101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101000101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101000101000101) && ({row_reg, col_reg}<19'b0011101000101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101000101010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101000101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011101000101010101) && ({row_reg, col_reg}<19'b0011101000101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101000101011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101000101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000101011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011101000101011100) && ({row_reg, col_reg}<19'b0011101000101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101000101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101000101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101000101100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101000101100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000101100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101000101100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101000101100111) && ({row_reg, col_reg}<19'b0011101000101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101000101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101000101101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101000101101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101000101101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011101000101101111) && ({row_reg, col_reg}<19'b0011101000101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101000101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101000101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000101111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101000101111010) && ({row_reg, col_reg}<19'b0011101000101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101000101111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000101111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011101000110000000) && ({row_reg, col_reg}<19'b0011101000110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101000110110000) && ({row_reg, col_reg}<19'b0011101000110110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011101000110110010) && ({row_reg, col_reg}<19'b0011101000110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101000110111000)) color_data = 12'b000100110011;
		if(({row_reg, col_reg}==19'b0011101000110111001)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}==19'b0011101000110111010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0011101000110111011) && ({row_reg, col_reg}<19'b0011101000110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101000110111110) && ({row_reg, col_reg}<19'b0011101000111000000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011101000111000000) && ({row_reg, col_reg}<19'b0011101001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101001001010001) && ({row_reg, col_reg}<19'b0011101001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011101001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011101001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011101010000000000) && ({row_reg, col_reg}<19'b0011101010010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101010010110001) && ({row_reg, col_reg}<19'b0011101010010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101010010110100) && ({row_reg, col_reg}<19'b0011101010010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101010010110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101010010111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010010111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101010010111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101010010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101010010111100) && ({row_reg, col_reg}<19'b0011101010011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010011000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101010011000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101010011000010) && ({row_reg, col_reg}<19'b0011101010011000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010011000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101010011000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011101010011000110) && ({row_reg, col_reg}<19'b0011101010011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101010011001111) && ({row_reg, col_reg}<19'b0011101010011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101010011010001) && ({row_reg, col_reg}<19'b0011101010011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101010011011010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101010011011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010011011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101010011011101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101010011011110) && ({row_reg, col_reg}<19'b0011101010011100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010011100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101010011100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101010011100010) && ({row_reg, col_reg}<19'b0011101010011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010011100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101010011100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101010011100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101010011100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101010011101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101010011101001) && ({row_reg, col_reg}<19'b0011101010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101010011111011) && ({row_reg, col_reg}<19'b0011101010011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010011111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010011111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010011111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101010100000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101010100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011101010100000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010100000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101010100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101010100000110) && ({row_reg, col_reg}<19'b0011101010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101010100010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101010100010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010100010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101010100010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101010100010111) && ({row_reg, col_reg}<19'b0011101010100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010100011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101010100011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011101010100011011) && ({row_reg, col_reg}<19'b0011101010100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101010100011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010100100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101010100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101010100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101010100100100) && ({row_reg, col_reg}<19'b0011101010100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101010100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101010100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101010100101011) && ({row_reg, col_reg}<19'b0011101010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101010100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101010100110001) && ({row_reg, col_reg}<19'b0011101010100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101010100110110) && ({row_reg, col_reg}<19'b0011101010100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101010100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011101010100111111) && ({row_reg, col_reg}<19'b0011101010101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010101000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101010101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101010101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101010101000101) && ({row_reg, col_reg}<19'b0011101010101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101010101010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101010101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011101010101010101) && ({row_reg, col_reg}<19'b0011101010101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010101011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101010101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010101011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011101010101011100) && ({row_reg, col_reg}<19'b0011101010101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101010101011111) && ({row_reg, col_reg}<19'b0011101010101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010101100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101010101100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101010101100011) && ({row_reg, col_reg}<19'b0011101010101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010101100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101010101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101010101100111) && ({row_reg, col_reg}<19'b0011101010101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010101101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101010101101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010101101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101010101101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011101010101101111) && ({row_reg, col_reg}<19'b0011101010101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101010101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101010101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011101010101111010) && ({row_reg, col_reg}<19'b0011101010101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101010101111101) && ({row_reg, col_reg}<19'b0011101010101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101010110000000) && ({row_reg, col_reg}<19'b0011101010110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101010110110000) && ({row_reg, col_reg}<19'b0011101010110110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011101010110110010) && ({row_reg, col_reg}<19'b0011101010110110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101010110110101) && ({row_reg, col_reg}<19'b0011101010110111000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011101010110111000)) color_data = 12'b001101010110;
		if(({row_reg, col_reg}==19'b0011101010110111001)) color_data = 12'b001001000101;
		if(({row_reg, col_reg}==19'b0011101010110111010)) color_data = 12'b000100100011;
		if(({row_reg, col_reg}==19'b0011101010110111011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011101010110111100) && ({row_reg, col_reg}<19'b0011101010110111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101010110111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0011101010111000000) && ({row_reg, col_reg}<19'b0011101011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101011001010001) && ({row_reg, col_reg}<19'b0011101011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011101011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011101011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011101100000000000) && ({row_reg, col_reg}<19'b0011101100010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101100010110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101100010111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101100010111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101100010111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101100010111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011101100010111100) && ({row_reg, col_reg}<19'b0011101100011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100011000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101100011000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101100011000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101100011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100011000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101100011000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101100011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100011000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101100011001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101100011001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101100011001010) && ({row_reg, col_reg}<19'b0011101100011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101100011001111) && ({row_reg, col_reg}<19'b0011101100011010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101100011010001) && ({row_reg, col_reg}<19'b0011101100011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100011010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101100011010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101100011011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011101100011011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101100011011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011101100011011011) && ({row_reg, col_reg}<19'b0011101100011011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100011011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101100011011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101100011011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101100011100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101100011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101100011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100011100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101100011100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101100011100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101100011100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101100011100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011101100011101000) && ({row_reg, col_reg}<19'b0011101100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100011101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101100011101110) && ({row_reg, col_reg}<19'b0011101100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101100011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101100011111010) && ({row_reg, col_reg}<19'b0011101100011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101100011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100011111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101100011111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101100011111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101100100000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100100000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101100100000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101100100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101100100000111) && ({row_reg, col_reg}<19'b0011101100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101100100010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100100010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101100100010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100100010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101100100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101100100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101100100011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101100100011010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101100100011011) && ({row_reg, col_reg}<19'b0011101100100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101100100011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101100100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100100100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011101100100100001) && ({row_reg, col_reg}<19'b0011101100100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101100100100100) && ({row_reg, col_reg}<19'b0011101100100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101100100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101100100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101100100101011) && ({row_reg, col_reg}<19'b0011101100100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101100100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101100100110001) && ({row_reg, col_reg}<19'b0011101100100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101100100110110) && ({row_reg, col_reg}<19'b0011101100100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101100100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011101100100111111) && ({row_reg, col_reg}<19'b0011101100101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100101000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101100101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101100101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101100101000101) && ({row_reg, col_reg}<19'b0011101100101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101100101010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011101100101010011) && ({row_reg, col_reg}<19'b0011101100101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101100101010110) && ({row_reg, col_reg}<19'b0011101100101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100101011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100101011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011101100101011100) && ({row_reg, col_reg}<19'b0011101100101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101100101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100101100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101100101100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100101100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101100101100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100101100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101100101100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011101100101100110) && ({row_reg, col_reg}<19'b0011101100101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101100101101001) && ({row_reg, col_reg}<19'b0011101100101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100101101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100101101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100101101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101100101101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101100101101111) && ({row_reg, col_reg}<19'b0011101100101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101100101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101100101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101100101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101100101111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101100101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101100101111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011101100101111101) && ({row_reg, col_reg}<19'b0011101100101111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011101100101111111) && ({row_reg, col_reg}<19'b0011101100110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101100110110011) && ({row_reg, col_reg}<19'b0011101100110110110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011101100110110110) && ({row_reg, col_reg}<19'b0011101100110111000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0011101100110111000)) color_data = 12'b010110001001;
		if(({row_reg, col_reg}==19'b0011101100110111001)) color_data = 12'b010001101000;
		if(({row_reg, col_reg}==19'b0011101100110111010)) color_data = 12'b001001000101;
		if(({row_reg, col_reg}==19'b0011101100110111011)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}>=19'b0011101100110111100) && ({row_reg, col_reg}<19'b0011101101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101101001010001) && ({row_reg, col_reg}<19'b0011101101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011101101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011101101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011101110000000000) && ({row_reg, col_reg}<19'b0011101110010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101110010110011) && ({row_reg, col_reg}<19'b0011101110010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101110010110101) && ({row_reg, col_reg}<19'b0011101110010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110010111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101110010111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101110010111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011101110010111100) && ({row_reg, col_reg}<19'b0011101110010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101110010111111) && ({row_reg, col_reg}<19'b0011101110011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101110011000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011101110011000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011101110011000100) && ({row_reg, col_reg}<19'b0011101110011001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110011001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101110011001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110011001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101110011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101110011001100) && ({row_reg, col_reg}<19'b0011101110011010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110011010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110011010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101110011010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110011010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011101110011011000) && ({row_reg, col_reg}<19'b0011101110011011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110011011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101110011011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011101110011011111) && ({row_reg, col_reg}<19'b0011101110011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110011100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101110011100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101110011100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101110011100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101110011100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101110011101000) && ({row_reg, col_reg}<19'b0011101110011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110011101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101110011101110) && ({row_reg, col_reg}<19'b0011101110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110011111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011101110011111001) && ({row_reg, col_reg}<19'b0011101110011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110011111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101110011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110011111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101110011111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110100000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101110100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101110100000011) && ({row_reg, col_reg}<19'b0011101110100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110100000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110100000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101110100000111) && ({row_reg, col_reg}<19'b0011101110100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101110100010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110100010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101110100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101110100010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101110100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110100011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011101110100011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101110100011010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101110100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110100011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011101110100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101110100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110100100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011101110100100001) && ({row_reg, col_reg}<19'b0011101110100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101110100100100) && ({row_reg, col_reg}<19'b0011101110100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101110100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101110100101011) && ({row_reg, col_reg}<19'b0011101110100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101110100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101110100110001) && ({row_reg, col_reg}<19'b0011101110100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101110100110110) && ({row_reg, col_reg}<19'b0011101110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101110100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011101110100111111) && ({row_reg, col_reg}<19'b0011101110101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110101000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011101110101000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101110101000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101110101000101) && ({row_reg, col_reg}<19'b0011101110101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110101010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101110101010011) && ({row_reg, col_reg}<19'b0011101110101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101110101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101110101010111) && ({row_reg, col_reg}<19'b0011101110101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110101011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110101011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101110101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101110101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110101100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101110101100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101110101100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110101100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101110101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011101110101100101) && ({row_reg, col_reg}<19'b0011101110101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110101100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101110101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101110101101001) && ({row_reg, col_reg}<19'b0011101110101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110101101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110101101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110101101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011101110101101111) && ({row_reg, col_reg}<19'b0011101110101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011101110101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011101110101111000) && ({row_reg, col_reg}<19'b0011101110101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110101111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011101110101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011101110101111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101110101111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011101110101111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101110101111111) && ({row_reg, col_reg}<19'b0011101110110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011101110110110011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011101110110110100) && ({row_reg, col_reg}<19'b0011101110110110110)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0011101110110110110) && ({row_reg, col_reg}<19'b0011101110110111000)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0011101110110111000)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==19'b0011101110110111001)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==19'b0011101110110111010)) color_data = 12'b001101010111;
		if(({row_reg, col_reg}==19'b0011101110110111011)) color_data = 12'b000100100100;
		if(({row_reg, col_reg}==19'b0011101110110111100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011101110110111101) && ({row_reg, col_reg}<19'b0011101111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011101111001010001) && ({row_reg, col_reg}<19'b0011101111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011101111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011101111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011110000000000000) && ({row_reg, col_reg}<19'b0011110000010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000010111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110000010111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011110000010111010) && ({row_reg, col_reg}<19'b0011110000010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000010111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110000010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110000010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110000010111111) && ({row_reg, col_reg}<19'b0011110000011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110000011000001) && ({row_reg, col_reg}<19'b0011110000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110000011000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110000011000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011110000011000110) && ({row_reg, col_reg}<19'b0011110000011001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000011001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110000011001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110000011001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110000011001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000011001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011110000011010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110000011010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110000011010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110000011010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110000011010100) && ({row_reg, col_reg}<19'b0011110000011010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011110000011010110) && ({row_reg, col_reg}<19'b0011110000011011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000011011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110000011011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110000011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011110000011011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110000011011101) && ({row_reg, col_reg}<19'b0011110000011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110000011100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110000011100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110000011100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110000011100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110000011100100) && ({row_reg, col_reg}<19'b0011110000011100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110000011100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011110000011100111) && ({row_reg, col_reg}<19'b0011110000011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110000011111100) && ({row_reg, col_reg}<19'b0011110000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000011111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011110000011111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000100000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110000100000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110000100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110000100000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000100000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110000100000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011110000100000111) && ({row_reg, col_reg}<19'b0011110000100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110000100001001) && ({row_reg, col_reg}<19'b0011110000100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110000100001011) && ({row_reg, col_reg}<19'b0011110000100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000100001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011110000100001111) && ({row_reg, col_reg}<19'b0011110000100010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000100010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110000100010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011110000100010011) && ({row_reg, col_reg}<19'b0011110000100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000100010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110000100010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110000100010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110000100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000100011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011110000100011010) && ({row_reg, col_reg}<19'b0011110000100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000100011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110000100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110000100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000100100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110000100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110000100100010) && ({row_reg, col_reg}<19'b0011110000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110000100101000) && ({row_reg, col_reg}<19'b0011110000100101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110000100101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110000100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110000100101100) && ({row_reg, col_reg}<19'b0011110000100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110000100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000100110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110000100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110000100110100) && ({row_reg, col_reg}<19'b0011110000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110000100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110000100111001) && ({row_reg, col_reg}<19'b0011110000100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000100111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011110000100111111) && ({row_reg, col_reg}<19'b0011110000101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000101000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110000101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000101000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110000101000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011110000101000101) && ({row_reg, col_reg}<19'b0011110000101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110000101001000) && ({row_reg, col_reg}<19'b0011110000101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000101010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110000101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000101010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011110000101010011) && ({row_reg, col_reg}<19'b0011110000101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000101010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011110000101010110) && ({row_reg, col_reg}<19'b0011110000101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000101011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110000101011010) && ({row_reg, col_reg}<19'b0011110000101011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000101011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110000101011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000101011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011110000101011111) && ({row_reg, col_reg}<19'b0011110000101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000101100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110000101100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110000101100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011110000101100100) && ({row_reg, col_reg}<19'b0011110000101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110000101101000) && ({row_reg, col_reg}<19'b0011110000101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000101101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000101101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000101101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110000101101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110000101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110000101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110000101110001) && ({row_reg, col_reg}<19'b0011110000101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110000101110011) && ({row_reg, col_reg}<19'b0011110000101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000101110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110000101110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011110000101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110000101111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110000101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000101111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110000101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110000101111111) && ({row_reg, col_reg}<19'b0011110000110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110000110110001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0011110000110110010)) color_data = 12'b000100010011;
		if(({row_reg, col_reg}==19'b0011110000110110011)) color_data = 12'b000000010011;
		if(({row_reg, col_reg}==19'b0011110000110110100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0011110000110110101)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0011110000110110110)) color_data = 12'b000100110111;
		if(({row_reg, col_reg}==19'b0011110000110110111)) color_data = 12'b001101101010;
		if(({row_reg, col_reg}==19'b0011110000110111000)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==19'b0011110000110111001)) color_data = 12'b001101101001;
		if(({row_reg, col_reg}==19'b0011110000110111010)) color_data = 12'b000100110110;
		if(({row_reg, col_reg}==19'b0011110000110111011)) color_data = 12'b000000010100;
		if(({row_reg, col_reg}>=19'b0011110000110111100) && ({row_reg, col_reg}<19'b0011110000110111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011110000110111110) && ({row_reg, col_reg}<19'b0011110001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110001001010001) && ({row_reg, col_reg}<19'b0011110001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011110001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011110001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011110010000000000) && ({row_reg, col_reg}<19'b0011110010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010010111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011110010010111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110010010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010010111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110010010111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110010010111111) && ({row_reg, col_reg}<19'b0011110010011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010011000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110010011000111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011110010011001000) && ({row_reg, col_reg}<19'b0011110010011001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110010011001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011110010011001011) && ({row_reg, col_reg}<19'b0011110010011010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010011010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011110010011010110) && ({row_reg, col_reg}<19'b0011110010011011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110010011011000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110010011011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110010011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110010011011011) && ({row_reg, col_reg}<19'b0011110010011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010011100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110010011100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011110010011100011) && ({row_reg, col_reg}<19'b0011110010011100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110010011100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110010011100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011110010011100111) && ({row_reg, col_reg}<19'b0011110010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110010011111001) && ({row_reg, col_reg}<19'b0011110010011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110010011111100) && ({row_reg, col_reg}<19'b0011110010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010011111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110010011111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110010100000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010100000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011110010100000100) && ({row_reg, col_reg}<19'b0011110010100000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010100000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110010100001000) && ({row_reg, col_reg}<19'b0011110010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110010100001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110010100001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110010100001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110010100001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010100010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110010100010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011110010100010010) && ({row_reg, col_reg}<19'b0011110010100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010100010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110010100010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110010100010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011110010100010111) && ({row_reg, col_reg}<19'b0011110010100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010100011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110010100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010100011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110010100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011110010100100000) && ({row_reg, col_reg}<19'b0011110010100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110010100100010) && ({row_reg, col_reg}<19'b0011110010100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110010100101000) && ({row_reg, col_reg}<19'b0011110010100101010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110010100101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110010100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110010100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110010100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110010100101111) && ({row_reg, col_reg}<19'b0011110010100110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110010100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110010100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110010100110100) && ({row_reg, col_reg}<19'b0011110010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110010100111001) && ({row_reg, col_reg}<19'b0011110010100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010100111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110010100111111) && ({row_reg, col_reg}<19'b0011110010101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010101000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110010101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010101000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110010101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110010101000101) && ({row_reg, col_reg}<19'b0011110010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010101010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011110010101010011) && ({row_reg, col_reg}<19'b0011110010101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010101010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011110010101010110) && ({row_reg, col_reg}<19'b0011110010101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010101011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110010101011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011110010101011011) && ({row_reg, col_reg}<19'b0011110010101100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010101100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110010101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110010101100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011110010101100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110010101100100) && ({row_reg, col_reg}<19'b0011110010101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010101100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110010101100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110010101101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011110010101101001) && ({row_reg, col_reg}<19'b0011110010101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010101101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110010101101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010101101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011110010101101110) && ({row_reg, col_reg}<19'b0011110010101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110010101110001) && ({row_reg, col_reg}<19'b0011110010101110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110010101110011) && ({row_reg, col_reg}<19'b0011110010101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010101110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110010101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110010101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010101111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110010101111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110010101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010101111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110010101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110010101111111) && ({row_reg, col_reg}<19'b0011110010110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110010110110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110010110110001)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0011110010110110010)) color_data = 12'b000100100011;
		if(({row_reg, col_reg}==19'b0011110010110110011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0011110010110110100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0011110010110110101)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0011110010110110110)) color_data = 12'b000100111000;
		if(({row_reg, col_reg}>=19'b0011110010110110111) && ({row_reg, col_reg}<19'b0011110010110111001)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==19'b0011110010110111001)) color_data = 12'b001101101010;
		if(({row_reg, col_reg}==19'b0011110010110111010)) color_data = 12'b000100110111;
		if(({row_reg, col_reg}==19'b0011110010110111011)) color_data = 12'b000000010100;
		if(({row_reg, col_reg}==19'b0011110010110111100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0011110010110111101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011110010110111110) && ({row_reg, col_reg}<19'b0011110011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110011001010001) && ({row_reg, col_reg}<19'b0011110011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011110011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011110011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011110100000000000) && ({row_reg, col_reg}<19'b0011110100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110100010111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100010111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110100010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100010111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110100010111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110100010111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011110100011000000) && ({row_reg, col_reg}<19'b0011110100011001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100011001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100011001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110100011001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011110100011001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110100011001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011110100011001101) && ({row_reg, col_reg}<19'b0011110100011001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100011001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110100011010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100011010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110100011010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110100011010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110100011010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100011010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011110100011010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110100011010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110100011011000) && ({row_reg, col_reg}<19'b0011110100011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100011100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011110100011100010) && ({row_reg, col_reg}<19'b0011110100011100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100011100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110100011100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011110100011100110) && ({row_reg, col_reg}<19'b0011110100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110100011111001) && ({row_reg, col_reg}<19'b0011110100011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110100011111011) && ({row_reg, col_reg}<19'b0011110100011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110100011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100011111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100011111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100100000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100100000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110100100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100100000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011110100100000101) && ({row_reg, col_reg}<19'b0011110100100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100100000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011110100100001000) && ({row_reg, col_reg}<19'b0011110100100001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100100001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110100100001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110100100001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110100100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100100001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110100100001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100100010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011110100100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110100100010010) && ({row_reg, col_reg}<19'b0011110100100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100100010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011110100100010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011110100100010110) && ({row_reg, col_reg}<19'b0011110100100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110100100011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100100011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110100100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100100011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011110100100011110) && ({row_reg, col_reg}<19'b0011110100100100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110100100100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110100100100010) && ({row_reg, col_reg}<19'b0011110100100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100100101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110100100101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110100100101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110100100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110100100101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100100110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110100100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110100100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110100100110100) && ({row_reg, col_reg}<19'b0011110100100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110100100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110100100111001) && ({row_reg, col_reg}<19'b0011110100100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100100111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110100100111111) && ({row_reg, col_reg}<19'b0011110100101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100101000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110100101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100101000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110100101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110100101000101) && ({row_reg, col_reg}<19'b0011110100101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100101010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110100101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011110100101010110) && ({row_reg, col_reg}<19'b0011110100101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110100101011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011110100101011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011110100101011100) && ({row_reg, col_reg}<19'b0011110100101011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110100101011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110100101011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110100101100000) && ({row_reg, col_reg}<19'b0011110100101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110100101100011) && ({row_reg, col_reg}<19'b0011110100101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100101100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110100101100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110100101101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100101101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110100101101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100101101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100101101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100101101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110100101110000) && ({row_reg, col_reg}<19'b0011110100101110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110100101110011) && ({row_reg, col_reg}<19'b0011110100101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110100101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110100101110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110100101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110100101111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110100101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110100101111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110100101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011110100101111111) && ({row_reg, col_reg}<19'b0011110100110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110100110110000) && ({row_reg, col_reg}<19'b0011110100110110010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0011110100110110010)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}==19'b0011110100110110011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0011110100110110100)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0011110100110110101)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==19'b0011110100110110110)) color_data = 12'b000100111001;
		if(({row_reg, col_reg}>=19'b0011110100110110111) && ({row_reg, col_reg}<19'b0011110100110111001)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==19'b0011110100110111001)) color_data = 12'b001101101100;
		if(({row_reg, col_reg}==19'b0011110100110111010)) color_data = 12'b001001001001;
		if(({row_reg, col_reg}==19'b0011110100110111011)) color_data = 12'b000000100110;
		if(({row_reg, col_reg}==19'b0011110100110111100)) color_data = 12'b000000010011;
		if(({row_reg, col_reg}==19'b0011110100110111101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0011110100110111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011110100110111111) && ({row_reg, col_reg}<19'b0011110101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110101001010001) && ({row_reg, col_reg}<19'b0011110101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011110101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011110101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011110110000000000) && ({row_reg, col_reg}<19'b0011110110010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110110010111011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011110110010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110110010111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011110110010111110) && ({row_reg, col_reg}<19'b0011110110011000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110011000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110011000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011110110011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110110011000011) && ({row_reg, col_reg}<19'b0011110110011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110011000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110110011000111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011110110011001000) && ({row_reg, col_reg}<19'b0011110110011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110011001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110110011001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110110011001101) && ({row_reg, col_reg}<19'b0011110110011010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011110110011010000) && ({row_reg, col_reg}<19'b0011110110011010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110110011010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110011010100) && ({row_reg, col_reg}<19'b0011110110011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110110011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110011011010) && ({row_reg, col_reg}<19'b0011110110011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110011100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110110011100001) && ({row_reg, col_reg}<19'b0011110110011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110011100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110110011100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011110110011100101) && ({row_reg, col_reg}<19'b0011110110011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110011100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110110011101000) && ({row_reg, col_reg}<19'b0011110110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110110011111001) && ({row_reg, col_reg}<19'b0011110110011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110011111101) && ({row_reg, col_reg}<19'b0011110110011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110110100000000) && ({row_reg, col_reg}<19'b0011110110100000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110110100000011) && ({row_reg, col_reg}<19'b0011110110100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110110100000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011110110100000110) && ({row_reg, col_reg}<19'b0011110110100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110100001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011110110100001011) && ({row_reg, col_reg}<19'b0011110110100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110100001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110110100001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110110100001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110110100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110110100010001) && ({row_reg, col_reg}<19'b0011110110100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110100010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110110100010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110110100010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110110100010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110110100010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110110100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110100011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011110110100011010) && ({row_reg, col_reg}<19'b0011110110100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110100011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110110100011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110110100011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011110110100100000) && ({row_reg, col_reg}<19'b0011110110100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110100100010) && ({row_reg, col_reg}<19'b0011110110100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110110100101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011110110100101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110110100101011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110110100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110110100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110110100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110100110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110110100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110110100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110100110100) && ({row_reg, col_reg}<19'b0011110110100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110100110111) && ({row_reg, col_reg}<19'b0011110110100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011110110100111111) && ({row_reg, col_reg}<19'b0011110110101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110101000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110110101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110101000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110110101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110101000101) && ({row_reg, col_reg}<19'b0011110110101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110101010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110110101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110101010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110110101010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110110101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110101011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110110101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110101011010) && ({row_reg, col_reg}<19'b0011110110101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110101011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011110110101011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110110101011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011110110101011111) && ({row_reg, col_reg}<19'b0011110110101100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110101100001) && ({row_reg, col_reg}<19'b0011110110101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110110101100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011110110101100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011110110101100111) && ({row_reg, col_reg}<19'b0011110110101101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011110110101101001) && ({row_reg, col_reg}<19'b0011110110101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011110110101101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110110101101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110101101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011110110101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110101110000) && ({row_reg, col_reg}<19'b0011110110101110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011110110101110011) && ({row_reg, col_reg}<19'b0011110110101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011110110101110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011110110101111000) && ({row_reg, col_reg}<19'b0011110110101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110101111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110110101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110110101111100) && ({row_reg, col_reg}<19'b0011110110101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011110110101111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011110110101111111) && ({row_reg, col_reg}<19'b0011110110110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011110110110110001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011110110110110010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0011110110110110011)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0011110110110110100)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0011110110110110101)) color_data = 12'b000000010111;
		if(({row_reg, col_reg}==19'b0011110110110110110)) color_data = 12'b000101001011;
		if(({row_reg, col_reg}==19'b0011110110110110111)) color_data = 12'b001101101101;
		if(({row_reg, col_reg}==19'b0011110110110111000)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==19'b0011110110110111001)) color_data = 12'b001101101101;
		if(({row_reg, col_reg}==19'b0011110110110111010)) color_data = 12'b010001101100;
		if(({row_reg, col_reg}==19'b0011110110110111011)) color_data = 12'b001101011010;
		if(({row_reg, col_reg}==19'b0011110110110111100)) color_data = 12'b001101000111;
		if(({row_reg, col_reg}==19'b0011110110110111101)) color_data = 12'b000100100100;
		if(({row_reg, col_reg}==19'b0011110110110111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011110110110111111) && ({row_reg, col_reg}<19'b0011110111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011110111001010001) && ({row_reg, col_reg}<19'b0011110111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011110111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011110111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011111000000000000) && ({row_reg, col_reg}<19'b0011111000010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000010111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111000010111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000010111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011111000010111111) && ({row_reg, col_reg}<19'b0011111000011000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000011000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111000011000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111000011000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111000011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111000011000101) && ({row_reg, col_reg}<19'b0011111000011001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111000011001000) && ({row_reg, col_reg}<19'b0011111000011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111000011001100) && ({row_reg, col_reg}<19'b0011111000011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111000011010000) && ({row_reg, col_reg}<19'b0011111000011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111000011011000) && ({row_reg, col_reg}<19'b0011111000011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000011011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000011011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111000011011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011111000011011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111000011011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011111000011100000) && ({row_reg, col_reg}<19'b0011111000011100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000011100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111000011100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011111000011100100) && ({row_reg, col_reg}<19'b0011111000011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000011100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111000011101000) && ({row_reg, col_reg}<19'b0011111000011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111000011111001) && ({row_reg, col_reg}<19'b0011111000011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111000011111101) && ({row_reg, col_reg}<19'b0011111000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000100000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111000100000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111000100000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111000100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111000100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111000100000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011111000100001000) && ({row_reg, col_reg}<19'b0011111000100001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000100001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111000100001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111000100001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111000100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111000100001111) && ({row_reg, col_reg}<19'b0011111000100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000100010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111000100010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000100010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111000100010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111000100010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000100011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011111000100011010) && ({row_reg, col_reg}<19'b0011111000100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000100011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111000100011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111000100011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000100011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011111000100100000) && ({row_reg, col_reg}<19'b0011111000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111000100101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111000100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111000100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000100101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111000100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000100110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111000100110100) && ({row_reg, col_reg}<19'b0011111000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111000100110111) && ({row_reg, col_reg}<19'b0011111000100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111000100111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111000100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000100111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000101000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111000101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000101000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011111000101000100) && ({row_reg, col_reg}<19'b0011111000101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111000101000111) && ({row_reg, col_reg}<19'b0011111000101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111000101010001) && ({row_reg, col_reg}<19'b0011111000101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000101010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111000101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111000101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000101010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111000101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000101011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111000101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111000101011010) && ({row_reg, col_reg}<19'b0011111000101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000101100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111000101100001) && ({row_reg, col_reg}<19'b0011111000101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000101100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111000101100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011111000101100110) && ({row_reg, col_reg}<19'b0011111000101101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000101101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111000101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000101101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111000101101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111000101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111000101110000) && ({row_reg, col_reg}<19'b0011111000101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111000101111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011111000101111001) && ({row_reg, col_reg}<19'b0011111000101111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000101111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111000101111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111000101111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111000101111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111000101111111) && ({row_reg, col_reg}<19'b0011111000110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111000110110001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011111000110110010)) color_data = 12'b000100100100;
		if(({row_reg, col_reg}==19'b0011111000110110011)) color_data = 12'b001000110111;
		if(({row_reg, col_reg}==19'b0011111000110110100)) color_data = 12'b001001001001;
		if(({row_reg, col_reg}==19'b0011111000110110101)) color_data = 12'b001101011100;
		if(({row_reg, col_reg}==19'b0011111000110110110)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==19'b0011111000110110111)) color_data = 12'b010001111111;
		if(({row_reg, col_reg}==19'b0011111000110111000)) color_data = 12'b001001011101;
		if(({row_reg, col_reg}==19'b0011111000110111001)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==19'b0011111000110111010)) color_data = 12'b010110001110;
		if(({row_reg, col_reg}==19'b0011111000110111011)) color_data = 12'b011010001101;
		if(({row_reg, col_reg}==19'b0011111000110111100)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==19'b0011111000110111101)) color_data = 12'b001101000110;
		if(({row_reg, col_reg}==19'b0011111000110111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011111000110111111) && ({row_reg, col_reg}<19'b0011111001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111001001010001) && ({row_reg, col_reg}<19'b0011111001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011111001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011111001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011111010000000000) && ({row_reg, col_reg}<19'b0011111010010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111010010111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111010011000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011111010011000001) && ({row_reg, col_reg}<19'b0011111010011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010011000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111010011000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111010011000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010011000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011111010011000111) && ({row_reg, col_reg}<19'b0011111010011001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111010011001010) && ({row_reg, col_reg}<19'b0011111010011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111010011001100) && ({row_reg, col_reg}<19'b0011111010011011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010011011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111010011011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111010011011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111010011011101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111010011011110) && ({row_reg, col_reg}<19'b0011111010011100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010011100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111010011100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111010011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111010011100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111010011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111010011100111) && ({row_reg, col_reg}<19'b0011111010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111010011111001) && ({row_reg, col_reg}<19'b0011111010100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010100000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011111010100000010) && ({row_reg, col_reg}<19'b0011111010100000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0011111010100000101) && ({row_reg, col_reg}<19'b0011111010100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111010100001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111010100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011111010100001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111010100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111010100001100) && ({row_reg, col_reg}<19'b0011111010100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010100010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111010100010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111010100010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010100010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111010100010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010100010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111010100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010100011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111010100011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111010100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111010100011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010100011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011111010100100000) && ({row_reg, col_reg}<19'b0011111010100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010100101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111010100101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111010100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010100101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111010100101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111010100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010100110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111010100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111010100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111010100110100) && ({row_reg, col_reg}<19'b0011111010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111010100110111) && ({row_reg, col_reg}<19'b0011111010100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111010100111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011111010100111101) && ({row_reg, col_reg}<19'b0011111010100111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011111010100111111) && ({row_reg, col_reg}<19'b0011111010101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111010101000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111010101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010101000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011111010101000100) && ({row_reg, col_reg}<19'b0011111010101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111010101000111) && ({row_reg, col_reg}<19'b0011111010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111010101010001) && ({row_reg, col_reg}<19'b0011111010101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010101010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111010101010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111010101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010101010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111010101010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011111010101011000) && ({row_reg, col_reg}<19'b0011111010101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111010101011100) && ({row_reg, col_reg}<19'b0011111010101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111010101011110) && ({row_reg, col_reg}<19'b0011111010101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111010101100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111010101100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011111010101100101) && ({row_reg, col_reg}<19'b0011111010101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010101101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111010101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010101101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111010101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010101101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111010101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111010101101110) && ({row_reg, col_reg}<19'b0011111010101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111010101110000) && ({row_reg, col_reg}<19'b0011111010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010101111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111010101111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111010101111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111010101111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111010101111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111010101111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111010101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111010110000000) && ({row_reg, col_reg}<19'b0011111010110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111010110110001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0011111010110110010)) color_data = 12'b001000110101;
		if(({row_reg, col_reg}==19'b0011111010110110011)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==19'b0011111010110110100)) color_data = 12'b011010001101;
		if(({row_reg, col_reg}==19'b0011111010110110101)) color_data = 12'b011010001111;
		if(({row_reg, col_reg}==19'b0011111010110110110)) color_data = 12'b010110001111;
		if(({row_reg, col_reg}==19'b0011111010110110111)) color_data = 12'b010001111111;
		if(({row_reg, col_reg}==19'b0011111010110111000)) color_data = 12'b001001011110;
		if(({row_reg, col_reg}==19'b0011111010110111001)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==19'b0011111010110111010)) color_data = 12'b010101111110;
		if(({row_reg, col_reg}==19'b0011111010110111011)) color_data = 12'b010101111101;
		if(({row_reg, col_reg}==19'b0011111010110111100)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==19'b0011111010110111101)) color_data = 12'b001000110101;
		if(({row_reg, col_reg}==19'b0011111010110111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011111010110111111) && ({row_reg, col_reg}<19'b0011111011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111011001010001) && ({row_reg, col_reg}<19'b0011111011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011111011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011111011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011111100000000000) && ({row_reg, col_reg}<19'b0011111100011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100011000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011111100011000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100011000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111100011000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011111100011000100) && ({row_reg, col_reg}<19'b0011111100011000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100011000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111100011000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0011111100011001000) && ({row_reg, col_reg}<19'b0011111100011001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0011111100011001010) && ({row_reg, col_reg}<19'b0011111100011001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011111100011001101) && ({row_reg, col_reg}<19'b0011111100011010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011111100011010000) && ({row_reg, col_reg}<19'b0011111100011010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111100011010011) && ({row_reg, col_reg}<19'b0011111100011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111100011010101) && ({row_reg, col_reg}<19'b0011111100011010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111100011010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111100011011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111100011011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111100011011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111100011011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111100011011100) && ({row_reg, col_reg}<19'b0011111100011011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100011011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111100011011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111100011100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111100011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111100011100010) && ({row_reg, col_reg}<19'b0011111100011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111100011100100) && ({row_reg, col_reg}<19'b0011111100011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111100011100110) && ({row_reg, col_reg}<19'b0011111100011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100100000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111100100000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111100100000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100100000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111100100000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0011111100100000110) && ({row_reg, col_reg}<19'b0011111100100001000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0011111100100001000) && ({row_reg, col_reg}<19'b0011111100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111100100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111100100010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111100100010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100100010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111100100010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100100010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111100100010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011111100100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111100100010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111100100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111100100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100100011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100100011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111100100011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111100100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111100100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011111100100011111) && ({row_reg, col_reg}<19'b0011111100100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100100101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111100100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100100101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111100100101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111100100101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111100100101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111100100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100100110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111100100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111100100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111100100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111100100110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111100100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111100100111001) && ({row_reg, col_reg}<19'b0011111100100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100100111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011111100100111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111100100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100100111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011111100101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111100101000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111100101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100101000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111100101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100101000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111100101000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111100101000111) && ({row_reg, col_reg}<19'b0011111100101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111100101010010) && ({row_reg, col_reg}<19'b0011111100101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100101010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011111100101010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111100101010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111100101010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111100101011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111100101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111100101011010) && ({row_reg, col_reg}<19'b0011111100101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111100101011100) && ({row_reg, col_reg}<19'b0011111100101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111100101011110) && ({row_reg, col_reg}<19'b0011111100101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100101100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111100101100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111100101100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0011111100101100100) && ({row_reg, col_reg}<19'b0011111100101100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111100101100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100101101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111100101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111100101101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111100101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100101101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111100101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100101101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011111100101101111) && ({row_reg, col_reg}<19'b0011111100101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100101111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111100101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100101111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111100101111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111100101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111100101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100101111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111100110000000) && ({row_reg, col_reg}<19'b0011111100110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111100110110001)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}==19'b0011111100110110010)) color_data = 12'b000100100101;
		if(({row_reg, col_reg}==19'b0011111100110110011)) color_data = 12'b001101001000;
		if(({row_reg, col_reg}==19'b0011111100110110100)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==19'b0011111100110110101)) color_data = 12'b010001101101;
		if(({row_reg, col_reg}==19'b0011111100110110110)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==19'b0011111100110110111)) color_data = 12'b001001011111;
		if(({row_reg, col_reg}==19'b0011111100110111000)) color_data = 12'b001101101111;
		if(({row_reg, col_reg}==19'b0011111100110111001)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==19'b0011111100110111010)) color_data = 12'b001001011100;
		if(({row_reg, col_reg}==19'b0011111100110111011)) color_data = 12'b001001001001;
		if(({row_reg, col_reg}==19'b0011111100110111100)) color_data = 12'b000100100110;
		if(({row_reg, col_reg}==19'b0011111100110111101)) color_data = 12'b000000010011;
		if(({row_reg, col_reg}==19'b0011111100110111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011111100110111111) && ({row_reg, col_reg}<19'b0011111101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111101001010001) && ({row_reg, col_reg}<19'b0011111101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011111101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011111101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0011111110000000000) && ({row_reg, col_reg}<19'b0011111110010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111110010111001) && ({row_reg, col_reg}<19'b0011111110010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111110010111110) && ({row_reg, col_reg}<19'b0011111110011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111110011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111110011000010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011111110011000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111110011000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111110011000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111110011000110) && ({row_reg, col_reg}<19'b0011111110011010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0011111110011010001) && ({row_reg, col_reg}<19'b0011111110011010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011111110011010101) && ({row_reg, col_reg}<19'b0011111110011011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110011011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111110011011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111110011011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111110011011111) && ({row_reg, col_reg}<19'b0011111110011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111110011100010) && ({row_reg, col_reg}<19'b0011111110011100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111110011100100) && ({row_reg, col_reg}<19'b0011111110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111110011111011) && ({row_reg, col_reg}<19'b0011111110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111110011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111110100000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011111110100000001) && ({row_reg, col_reg}<19'b0011111110100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111110100000100) && ({row_reg, col_reg}<19'b0011111110100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110100000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111110100001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111110100001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111110100001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111110100001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110100001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111110100001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111110100001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111110100001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110100010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111110100010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111110100010010) && ({row_reg, col_reg}<19'b0011111110100010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110100010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111110100010101) && ({row_reg, col_reg}<19'b0011111110100010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110100010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111110100011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111110100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110100011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111110100011011) && ({row_reg, col_reg}<19'b0011111110100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111110100011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0011111110100011111) && ({row_reg, col_reg}<19'b0011111110100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110100101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111110100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110100101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111110100101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111110100101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111110100101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110100101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111110100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111110100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111110100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0011111110100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111110100110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111110100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111110100111001) && ({row_reg, col_reg}<19'b0011111110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110100111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111110100111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111110100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110100111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0011111110101000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111110101000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0011111110101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110101000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0011111110101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110101000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111110101000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111110101000111) && ({row_reg, col_reg}<19'b0011111110101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111110101010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0011111110101010011) && ({row_reg, col_reg}<19'b0011111110101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110101010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0011111110101010111) && ({row_reg, col_reg}<19'b0011111110101011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110101011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111110101011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011111110101011011) && ({row_reg, col_reg}<19'b0011111110101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111110101011110) && ({row_reg, col_reg}<19'b0011111110101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110101100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0011111110101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111110101100010) && ({row_reg, col_reg}<19'b0011111110101100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110101100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111110101100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111110101100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111110101100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111110101101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111110101101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0011111110101101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0011111110101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110101101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0011111110101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110101101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0011111110101101111) && ({row_reg, col_reg}<19'b0011111110101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111110101111010) && ({row_reg, col_reg}<19'b0011111110101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0011111110101111101) && ({row_reg, col_reg}<19'b0011111110101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110101111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0011111110110000000) && ({row_reg, col_reg}<19'b0011111110110110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0011111110110110010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0011111110110110011)) color_data = 12'b000000010100;
		if(({row_reg, col_reg}==19'b0011111110110110100)) color_data = 12'b000000100110;
		if(({row_reg, col_reg}==19'b0011111110110110101)) color_data = 12'b000100101000;
		if(({row_reg, col_reg}>=19'b0011111110110110110) && ({row_reg, col_reg}<19'b0011111110110111000)) color_data = 12'b000000101001;
		if(({row_reg, col_reg}==19'b0011111110110111000)) color_data = 12'b010101111110;
		if(({row_reg, col_reg}==19'b0011111110110111001)) color_data = 12'b001101011100;
		if(({row_reg, col_reg}==19'b0011111110110111010)) color_data = 12'b000100111000;
		if(({row_reg, col_reg}==19'b0011111110110111011)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==19'b0011111110110111100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0011111110110111101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0011111110110111110) && ({row_reg, col_reg}<19'b0011111111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0011111111001010001) && ({row_reg, col_reg}<19'b0011111111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0011111111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0011111111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100000000000000000) && ({row_reg, col_reg}<19'b0100000000011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000000011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000000011000001) && ({row_reg, col_reg}<19'b0100000000011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000000011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000000011000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100000000011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000011000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000000011001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0100000000011001001) && ({row_reg, col_reg}<19'b0100000000011001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000000011001100) && ({row_reg, col_reg}<19'b0100000000011001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0100000000011001110) && ({row_reg, col_reg}<19'b0100000000011011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000011011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000000011011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000000011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000000011011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100000000011011101) && ({row_reg, col_reg}<19'b0100000000011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000000011100000) && ({row_reg, col_reg}<19'b0100000000100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000000100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000000100000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000000100000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000000100000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100000000100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000100001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0100000000100001001) && ({row_reg, col_reg}<19'b0100000000100001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000100001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100000000100010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000100010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100000000100010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000000100010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000000100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000000100010101) && ({row_reg, col_reg}<19'b0100000000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000000100011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100000000100011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000000100011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000000100011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000000100011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000000100011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000000100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000000100011111) && ({row_reg, col_reg}<19'b0100000000100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000000100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000000100101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100000000100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000000100101100) && ({row_reg, col_reg}<19'b0100000000100101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000100101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000000100101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0100000000100110000) && ({row_reg, col_reg}<19'b0100000000100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000000100111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000000100111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000000100111111) && ({row_reg, col_reg}<19'b0100000000101000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000101000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100000000101000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000000101000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100000000101000100) && ({row_reg, col_reg}<19'b0100000000101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000000101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000000101000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100000000101001000) && ({row_reg, col_reg}<19'b0100000000101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000000101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000000101010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000101010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0100000000101011000) && ({row_reg, col_reg}<19'b0100000000101011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0100000000101011011) && ({row_reg, col_reg}<19'b0100000000101011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0100000000101011101) && ({row_reg, col_reg}<19'b0100000000101011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100000000101011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0100000000101100000) && ({row_reg, col_reg}<19'b0100000000101100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000101100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100000000101100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100000000101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000000101100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000000101100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000101101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000000101101001) && ({row_reg, col_reg}<19'b0100000000101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000101101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000000101101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100000000101101101) && ({row_reg, col_reg}<19'b0100000000110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000000110110011) && ({row_reg, col_reg}<19'b0100000000110110101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0100000000110110101) && ({row_reg, col_reg}<19'b0100000000110111000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0100000000110111000)) color_data = 12'b000100100100;
		if(({row_reg, col_reg}>=19'b0100000000110111001) && ({row_reg, col_reg}<19'b0100000000110111011)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==19'b0100000000110111011)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==19'b0100000000110111100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100000000110111101)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0100000000110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000000110111111) && ({row_reg, col_reg}<19'b0100000001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000001001010001) && ({row_reg, col_reg}<19'b0100000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100000001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100000001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100000010000000000) && ({row_reg, col_reg}<19'b0100000010011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000010011000000) && ({row_reg, col_reg}<19'b0100000010011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000010011000010) && ({row_reg, col_reg}<19'b0100000010011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000010011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000010011000111) && ({row_reg, col_reg}<19'b0100000010011001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100000010011001011) && ({row_reg, col_reg}<19'b0100000010011001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100000010011001101) && ({row_reg, col_reg}<19'b0100000010011010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100000010011010000) && ({row_reg, col_reg}<19'b0100000010011011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000010011011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100000010011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000010011011011) && ({row_reg, col_reg}<19'b0100000010100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000010100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000010100000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100000010100000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100000010100001000) && ({row_reg, col_reg}<19'b0100000010100001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0100000010100001011) && ({row_reg, col_reg}<19'b0100000010100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000010100001101) && ({row_reg, col_reg}<19'b0100000010100010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000010100010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100000010100010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000010100010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100000010100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000010100010100) && ({row_reg, col_reg}<19'b0100000010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000010100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000010100011011) && ({row_reg, col_reg}<19'b0100000010100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000010100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000010100011110) && ({row_reg, col_reg}<19'b0100000010100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000010100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000010100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100000010100101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000010100101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000010100101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100000010100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100000010100110000) && ({row_reg, col_reg}<19'b0100000010100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000010100111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100000010100111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0100000010100111111) && ({row_reg, col_reg}<19'b0100000010101000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000010101000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100000010101000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010101000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100000010101000100) && ({row_reg, col_reg}<19'b0100000010101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000010101000110) && ({row_reg, col_reg}<19'b0100000010101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000010101001000) && ({row_reg, col_reg}<19'b0100000010101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000010101010001) && ({row_reg, col_reg}<19'b0100000010101010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000010101010011) && ({row_reg, col_reg}<19'b0100000010101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000010101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000010101010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100000010101011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000010101011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000010101011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000010101011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0100000010101011100) && ({row_reg, col_reg}<19'b0100000010101011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000010101011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100000010101011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100000010101100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000010101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000010101100010) && ({row_reg, col_reg}<19'b0100000010101100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000010101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000010101100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100000010101100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0100000010101101000) && ({row_reg, col_reg}<19'b0100000010101101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000010101101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100000010101101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000010101101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100000010101101101) && ({row_reg, col_reg}<19'b0100000010110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000010110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000010110111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100000010110111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010110111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100000010110111100) && ({row_reg, col_reg}<19'b0100000010110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000010110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000010110111111) && ({row_reg, col_reg}<19'b0100000011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000011001010001) && ({row_reg, col_reg}<19'b0100000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100000011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100000011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100000100000000000) && ({row_reg, col_reg}<19'b0100000100011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000100011000000) && ({row_reg, col_reg}<19'b0100000100011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100011000010) && ({row_reg, col_reg}<19'b0100000100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000100100000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000100100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100100000010) && ({row_reg, col_reg}<19'b0100000100100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000100100010110) && ({row_reg, col_reg}<19'b0100000100100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100100011000) && ({row_reg, col_reg}<19'b0100000100100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000100100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000100100011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100000100100100000) && ({row_reg, col_reg}<19'b0100000100100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000100100101100) && ({row_reg, col_reg}<19'b0100000100100101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000100100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100100101111) && ({row_reg, col_reg}<19'b0100000100100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000100100111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000100100111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100000100100111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000100101000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000100101000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000100101000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100000100101000011) && ({row_reg, col_reg}<19'b0100000100101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100101000110) && ({row_reg, col_reg}<19'b0100000100101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000100101010010) && ({row_reg, col_reg}<19'b0100000100101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100101010100) && ({row_reg, col_reg}<19'b0100000100101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000100101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000100101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000100101011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000100101011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000100101011100) && ({row_reg, col_reg}<19'b0100000100101011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000100101011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000100101011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000100101100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000100101100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000100101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000100101100011) && ({row_reg, col_reg}<19'b0100000100101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000100101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000100101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000100101100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100000100101101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000100101101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000100101101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000100101101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100000100101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100101101101) && ({row_reg, col_reg}<19'b0100000100101101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000100101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100101110000) && ({row_reg, col_reg}<19'b0100000100110111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000100110111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100000100110111010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100000100110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100110111100) && ({row_reg, col_reg}<19'b0100000100110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000100110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000100110111111) && ({row_reg, col_reg}<19'b0100000101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000101001010001) && ({row_reg, col_reg}<19'b0100000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100000101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100000101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100000110000000000) && ({row_reg, col_reg}<19'b0100000110011001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000110011001101) && ({row_reg, col_reg}<19'b0100000110011010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110011010000) && ({row_reg, col_reg}<19'b0100000110011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000110011011000) && ({row_reg, col_reg}<19'b0100000110011011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110011011110) && ({row_reg, col_reg}<19'b0100000110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000110100000000) && ({row_reg, col_reg}<19'b0100000110100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110100000101) && ({row_reg, col_reg}<19'b0100000110100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000110100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000110100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110100011010) && ({row_reg, col_reg}<19'b0100000110100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000110100011110) && ({row_reg, col_reg}<19'b0100000110100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110100100000) && ({row_reg, col_reg}<19'b0100000110100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000110100101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100000110100101001) && ({row_reg, col_reg}<19'b0100000110100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000110100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000110100111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100000110101000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100000110101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110101000010) && ({row_reg, col_reg}<19'b0100000110101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000110101000101) && ({row_reg, col_reg}<19'b0100000110101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110101000111) && ({row_reg, col_reg}<19'b0100000110101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000110101011011) && ({row_reg, col_reg}<19'b0100000110101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110101011110) && ({row_reg, col_reg}<19'b0100000110101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000110101100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100000110101100001) && ({row_reg, col_reg}<19'b0100000110101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000110101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110101100101) && ({row_reg, col_reg}<19'b0100000110101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000110101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100000110101101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100000110101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100000110101101010) && ({row_reg, col_reg}<19'b0100000110101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000110101101110) && ({row_reg, col_reg}<19'b0100000110101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110101110000) && ({row_reg, col_reg}<19'b0100000110110111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000110110111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100000110110111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100000110110111011) && ({row_reg, col_reg}<19'b0100000110110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100000110110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100000110110111111) && ({row_reg, col_reg}<19'b0100000111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100000111001010001) && ({row_reg, col_reg}<19'b0100000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100000111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100000111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100001000000000000) && ({row_reg, col_reg}<19'b0100001000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001000011000011) && ({row_reg, col_reg}<19'b0100001000011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000011001000) && ({row_reg, col_reg}<19'b0100001000100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001000100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000100001001) && ({row_reg, col_reg}<19'b0100001000100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100001000100001111) && ({row_reg, col_reg}<19'b0100001000100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000100010101) && ({row_reg, col_reg}<19'b0100001000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001000100011000) && ({row_reg, col_reg}<19'b0100001000100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000100011010) && ({row_reg, col_reg}<19'b0100001000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001000100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000100101001) && ({row_reg, col_reg}<19'b0100001000101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001000101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000101001000) && ({row_reg, col_reg}<19'b0100001000101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001000101010101) && ({row_reg, col_reg}<19'b0100001000101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000101011001) && ({row_reg, col_reg}<19'b0100001000101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001000101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000101101000) && ({row_reg, col_reg}<19'b0100001000101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001000101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000101101110) && ({row_reg, col_reg}<19'b0100001000110111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001000110111001) && ({row_reg, col_reg}<19'b0100001000110111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001000110111011) && ({row_reg, col_reg}<19'b0100001001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001001001010001) && ({row_reg, col_reg}<19'b0100001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100001001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100001001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100001010000000000) && ({row_reg, col_reg}<19'b0100001010100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001010100011011) && ({row_reg, col_reg}<19'b0100001010100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001010100011101) && ({row_reg, col_reg}<19'b0100001010101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001010101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100001010101000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100001010101000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100001010101000100) && ({row_reg, col_reg}<19'b0100001010101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001010101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001010101001000) && ({row_reg, col_reg}<19'b0100001010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001010101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100001010101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001010101010010) && ({row_reg, col_reg}<19'b0100001010101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001010101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001010101011001) && ({row_reg, col_reg}<19'b0100001010101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001010101011110) && ({row_reg, col_reg}<19'b0100001010101100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001010101100000) && ({row_reg, col_reg}<19'b0100001010101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001010101101011) && ({row_reg, col_reg}<19'b0100001010101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001010101101110) && ({row_reg, col_reg}<19'b0100001011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001011001010001) && ({row_reg, col_reg}<19'b0100001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100001011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100001011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100001100000000000) && ({row_reg, col_reg}<19'b0100001100011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001100011011100) && ({row_reg, col_reg}<19'b0100001100011011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001100011011110) && ({row_reg, col_reg}<19'b0100001100011100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100001100011100000) && ({row_reg, col_reg}<19'b0100001100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001100100000000) && ({row_reg, col_reg}<19'b0100001100100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001100100000100) && ({row_reg, col_reg}<19'b0100001100100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001100100001001) && ({row_reg, col_reg}<19'b0100001100100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001100100001111) && ({row_reg, col_reg}<19'b0100001100100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001100100011011) && ({row_reg, col_reg}<19'b0100001100100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001100100100000) && ({row_reg, col_reg}<19'b0100001100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001100101000000) && ({row_reg, col_reg}<19'b0100001100101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100001100101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100001100101000011) && ({row_reg, col_reg}<19'b0100001100101000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001100101000101) && ({row_reg, col_reg}<19'b0100001100101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001100101010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100001100101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001100101010010) && ({row_reg, col_reg}<19'b0100001100101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001100101100000) && ({row_reg, col_reg}<19'b0100001100101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001100101100010) && ({row_reg, col_reg}<19'b0100001100101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001100101101000) && ({row_reg, col_reg}<19'b0100001100101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001100101101011) && ({row_reg, col_reg}<19'b0100001100110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001100110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001100110111001) && ({row_reg, col_reg}<19'b0100001101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001101001010001) && ({row_reg, col_reg}<19'b0100001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100001101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100001101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100001110000000000) && ({row_reg, col_reg}<19'b0100001110011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001110011000110) && ({row_reg, col_reg}<19'b0100001110011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001110011001100) && ({row_reg, col_reg}<19'b0100001110100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001110100010000) && ({row_reg, col_reg}<19'b0100001110100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001110100010010) && ({row_reg, col_reg}<19'b0100001110100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001110100101000) && ({row_reg, col_reg}<19'b0100001110100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001110100101011) && ({row_reg, col_reg}<19'b0100001110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001110100111100) && ({row_reg, col_reg}<19'b0100001110100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001110100111110) && ({row_reg, col_reg}<19'b0100001110101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001110101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100001110101000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100001110101000110) && ({row_reg, col_reg}<19'b0100001110101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001110101010100) && ({row_reg, col_reg}<19'b0100001110101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001110101010110) && ({row_reg, col_reg}<19'b0100001110101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001110101011001) && ({row_reg, col_reg}<19'b0100001110101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001110101011100) && ({row_reg, col_reg}<19'b0100001110101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001110101100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100001110101100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001110101100010) && ({row_reg, col_reg}<19'b0100001110101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001110101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100001110101100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100001110101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100001110101100111) && ({row_reg, col_reg}<19'b0100001110101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100001110101101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100001110101110000) && ({row_reg, col_reg}<19'b0100001110110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001110110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001110110111001) && ({row_reg, col_reg}<19'b0100001110110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100001110110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100001110110111101) && ({row_reg, col_reg}<19'b0100001111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100001111001010001) && ({row_reg, col_reg}<19'b0100001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100001111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100001111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100010000000000000) && ({row_reg, col_reg}<19'b0100010000011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010000011110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100010000011111000) && ({row_reg, col_reg}<19'b0100010000011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010000011111101) && ({row_reg, col_reg}<19'b0100010000011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100010000011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010000100000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100010000100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010000100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100010000100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100010000100000100) && ({row_reg, col_reg}<19'b0100010000100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010000100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010000100000111) && ({row_reg, col_reg}<19'b0100010000100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010000100001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100010000100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100010000100001101) && ({row_reg, col_reg}<19'b0100010000100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010000100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100010000100010000) && ({row_reg, col_reg}<19'b0100010001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010001001010001) && ({row_reg, col_reg}<19'b0100010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100010001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100010001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100010010000000000) && ({row_reg, col_reg}<19'b0100010010011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010010011110011) && ({row_reg, col_reg}<19'b0100010010011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010010011110101) && ({row_reg, col_reg}<19'b0100010010011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010010011111001) && ({row_reg, col_reg}<19'b0100010010011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010010011111011) && ({row_reg, col_reg}<19'b0100010010011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010010011111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100010010011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100010010011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010010100000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100010010100000001) && ({row_reg, col_reg}<19'b0100010010100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010010100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010010100000100) && ({row_reg, col_reg}<19'b0100010010100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010010100000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100010010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100010010100001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100010010100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010010100001010) && ({row_reg, col_reg}<19'b0100010010100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010010100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010010100010000) && ({row_reg, col_reg}<19'b0100010011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010011001010001) && ({row_reg, col_reg}<19'b0100010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100010011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100010011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100010100000000000) && ({row_reg, col_reg}<19'b0100010100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010100011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010100011110001) && ({row_reg, col_reg}<19'b0100010100011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010100011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100010100011111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100010100011111011) && ({row_reg, col_reg}<19'b0100010100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010100100000001) && ({row_reg, col_reg}<19'b0100010100100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010100100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100010100100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010100100000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010100100001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100010100100001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010100100001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100010100100001011) && ({row_reg, col_reg}<19'b0100010101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010101001010001) && ({row_reg, col_reg}<19'b0100010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100010101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100010101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100010110000000000) && ({row_reg, col_reg}<19'b0100010110011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010110011110101) && ({row_reg, col_reg}<19'b0100010110011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010110011110111) && ({row_reg, col_reg}<19'b0100010110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010110011111010) && ({row_reg, col_reg}<19'b0100010110011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010110011111100) && ({row_reg, col_reg}<19'b0100010110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010110100000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100010110100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010110100000010) && ({row_reg, col_reg}<19'b0100010110100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100010110100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010110100000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100010110100000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0100010110100000111) && ({row_reg, col_reg}<19'b0100010110100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010110100001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100010110100001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100010110100001100) && ({row_reg, col_reg}<19'b0100010110100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100010110100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100010110100001111) && ({row_reg, col_reg}<19'b0100010111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100010111001010001) && ({row_reg, col_reg}<19'b0100010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100010111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100010111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100011000000000000) && ({row_reg, col_reg}<19'b0100011000011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011000011110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100011000011110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100011000011110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011000011110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011000011110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011000011110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100011000011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100011000011111000) && ({row_reg, col_reg}<19'b0100011000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011000100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100011000100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100011000100000010) && ({row_reg, col_reg}<19'b0100011000100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100011000100000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100011000100000110) && ({row_reg, col_reg}<19'b0100011000100001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011000100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0100011000100001001) && ({row_reg, col_reg}<19'b0100011000100001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011000100001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100011000100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011000100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100011000100001111) && ({row_reg, col_reg}<19'b0100011001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100011001001010001) && ({row_reg, col_reg}<19'b0100011001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100011001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100011001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100011010000000000) && ({row_reg, col_reg}<19'b0100011010011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011010011110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100011010011110010) && ({row_reg, col_reg}<19'b0100011010011110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011010011110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011010011110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100011010011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100011010011111001) && ({row_reg, col_reg}<19'b0100011010100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011010100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100011010100000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011010100000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011010100000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011010100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011010100001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011010100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011010100001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011010100001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100011010100001101) && ({row_reg, col_reg}<19'b0100011010100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011010100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100011010100010000) && ({row_reg, col_reg}<19'b0100011011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100011011001010001) && ({row_reg, col_reg}<19'b0100011011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100011011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100011011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100011100000000000) && ({row_reg, col_reg}<19'b0100011100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011100011110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100011100011110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011100011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011100011110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100011100011110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011100011110101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100011100011110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100011100011110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011100011111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100011100011111010) && ({row_reg, col_reg}<19'b0100011100011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011100011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100011100011111101) && ({row_reg, col_reg}<19'b0100011100100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011100100000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100011100100000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011100100000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011100100000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011100100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100011100100001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011100100001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011100100001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011100100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100011100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011100100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100011100100010000) && ({row_reg, col_reg}<19'b0100011101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100011101001010001) && ({row_reg, col_reg}<19'b0100011101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100011101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100011101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100011110000000000) && ({row_reg, col_reg}<19'b0100011110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011110011110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011110011110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100011110011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011110011110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100011110011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011110011110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100011110011110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100011110011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011110011111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011110011111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100011110011111010) && ({row_reg, col_reg}<19'b0100011110011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011110011111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100011110011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100011110011111110) && ({row_reg, col_reg}<19'b0100011110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011110100000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100011110100000001) && ({row_reg, col_reg}<19'b0100011110100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011110100000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100011110100000101) && ({row_reg, col_reg}<19'b0100011110100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011110100000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100011110100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100011110100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100011110100001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011110100001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011110100001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011110100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100011110100001110) && ({row_reg, col_reg}<19'b0100011111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100011111001010001) && ({row_reg, col_reg}<19'b0100011111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100011111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100011111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100100000000000000) && ({row_reg, col_reg}<19'b0100100000011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100000011101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100100000011101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100100000011110000) && ({row_reg, col_reg}<19'b0100100000011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100000011110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100100000011110011) && ({row_reg, col_reg}<19'b0100100000011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100000011110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100100000011110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100000011111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100100000011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100100000011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100000011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100000011111100) && ({row_reg, col_reg}<19'b0100100000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100000011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100000011111111) && ({row_reg, col_reg}<19'b0100100000100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100000100000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100100000100000101) && ({row_reg, col_reg}<19'b0100100000100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100000100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100100000100001000) && ({row_reg, col_reg}<19'b0100100000100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100000100001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000100001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100000100001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100100000100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100100000100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100000100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100100000100010000) && ({row_reg, col_reg}<19'b0100100001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100100001001010001) && ({row_reg, col_reg}<19'b0100100001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100100001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100100001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100100010000000000) && ({row_reg, col_reg}<19'b0100100010011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100010011101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100100010011101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100100010011110000) && ({row_reg, col_reg}<19'b0100100010011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100010011110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100100010011110011) && ({row_reg, col_reg}<19'b0100100010011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100010011110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100100010011110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100010011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100010011111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100100010011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100100010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100010011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100010011111100) && ({row_reg, col_reg}<19'b0100100010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100010011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100010011111111) && ({row_reg, col_reg}<19'b0100100010100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100010100000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100100010100000101) && ({row_reg, col_reg}<19'b0100100010100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100010100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100010100001000) && ({row_reg, col_reg}<19'b0100100010100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100010100001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100100010100001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100100010100001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100100010100001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100100010100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100010100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100010100010000) && ({row_reg, col_reg}<19'b0100100011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100100011001010001) && ({row_reg, col_reg}<19'b0100100011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100100011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100100011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100100100000000000) && ({row_reg, col_reg}<19'b0100100100011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100100011101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100100100011101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100100100011110000) && ({row_reg, col_reg}<19'b0100100100011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100100011110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100100100011110011) && ({row_reg, col_reg}<19'b0100100100011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100100011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100100100011110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100100100011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100100011111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100100100011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100100100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100100011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100100011111100) && ({row_reg, col_reg}<19'b0100100100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100100011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100100011111111) && ({row_reg, col_reg}<19'b0100100100100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100100100000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100100100100000101) && ({row_reg, col_reg}<19'b0100100100100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100100100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100100100001000) && ({row_reg, col_reg}<19'b0100100100100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100100100001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100100100100001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100100100100001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100100100100001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100100100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100100100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100100100010000) && ({row_reg, col_reg}<19'b0100100101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100100101001010001) && ({row_reg, col_reg}<19'b0100100101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100100101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100100101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100100110000000000) && ({row_reg, col_reg}<19'b0100100110011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100110011101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100100110011101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100100110011110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100110011110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100100110011110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0100100110011110011) && ({row_reg, col_reg}<19'b0100100110011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100110011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100100110011110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100100110011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100110011111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100100110011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100100110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100110011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100110011111100) && ({row_reg, col_reg}<19'b0100100110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100110011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100110011111111) && ({row_reg, col_reg}<19'b0100100110100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100110100000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100100110100000101) && ({row_reg, col_reg}<19'b0100100110100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100110100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100110100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100100110100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100100110100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100100110100001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100100110100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100110100001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100110100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100100110100001111) && ({row_reg, col_reg}<19'b0100100111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100100111001010001) && ({row_reg, col_reg}<19'b0100100111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100100111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100100111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100101000000000000) && ({row_reg, col_reg}<19'b0100101000011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101000011101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101000011101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100101000011110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101000011110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100101000011110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100101000011110011) && ({row_reg, col_reg}<19'b0100101000011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101000011110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100101000011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101000011111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100101000011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100101000011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101000011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101000011111100) && ({row_reg, col_reg}<19'b0100101000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101000011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101000011111111) && ({row_reg, col_reg}<19'b0100101000100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101000100000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100101000100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101000100000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100101000100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101000100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101000100001001) && ({row_reg, col_reg}<19'b0100101000100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101000100001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101000100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101000100001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101000100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100101000100001111) && ({row_reg, col_reg}<19'b0100101001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100101001001010001) && ({row_reg, col_reg}<19'b0100101001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100101001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100101001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100101010000000000) && ({row_reg, col_reg}<19'b0100101010011001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101010011001000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0100101010011001001) && ({row_reg, col_reg}<19'b0100101010011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101010011101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100101010011101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100101010011110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101010011110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100101010011110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100101010011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101010011110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101010011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101010011110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100101010011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101010011111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100101010011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100101010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101010011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101010011111100) && ({row_reg, col_reg}<19'b0100101010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101010011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101010011111111) && ({row_reg, col_reg}<19'b0100101010100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100101010100000010) && ({row_reg, col_reg}<19'b0100101010100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101010100000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100101010100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101010100000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100101010100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101010100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101010100001001) && ({row_reg, col_reg}<19'b0100101010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101010100001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101010100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101010100001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101010100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100101010100001111) && ({row_reg, col_reg}<19'b0100101011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100101011001010001) && ({row_reg, col_reg}<19'b0100101011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100101011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100101011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100101100000000000) && ({row_reg, col_reg}<19'b0100101100011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100101100011000101) && ({row_reg, col_reg}<19'b0100101100011001011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0100101100011001011) && ({row_reg, col_reg}<19'b0100101100011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101100011101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100101100011101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100101100011110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101100011110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101100011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100101100011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101100011110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101100011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101100011110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100101100011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101100011111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100101100011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100101100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101100011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101100011111100) && ({row_reg, col_reg}<19'b0100101100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101100011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101100011111111) && ({row_reg, col_reg}<19'b0100101100100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100101100100000010) && ({row_reg, col_reg}<19'b0100101100100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101100100000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100101100100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101100100000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100101100100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101100100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101100100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101100100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101100100001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101100100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101100100001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101100100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101100100001111) && ({row_reg, col_reg}<19'b0100101101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100101101001010001) && ({row_reg, col_reg}<19'b0100101101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100101101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100101101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100101110000000000) && ({row_reg, col_reg}<19'b0100101110011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100101110011000100) && ({row_reg, col_reg}<19'b0100101110011000110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0100101110011000110) && ({row_reg, col_reg}<19'b0100101110011001010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0100101110011001010) && ({row_reg, col_reg}<19'b0100101110011001100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0100101110011001100) && ({row_reg, col_reg}<19'b0100101110011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101110011101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100101110011101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100101110011110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101110011110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101110011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100101110011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101110011110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101110011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101110011110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100101110011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101110011111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100101110011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100101110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101110011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101110011111100) && ({row_reg, col_reg}<19'b0100101110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101110011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101110011111111) && ({row_reg, col_reg}<19'b0100101110100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100101110100000010) && ({row_reg, col_reg}<19'b0100101110100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101110100000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100101110100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101110100000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100101110100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101110100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100101110100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100101110100001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100101110100001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101110100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101110100001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101110100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100101110100001111) && ({row_reg, col_reg}<19'b0100101111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100101111001010001) && ({row_reg, col_reg}<19'b0100101111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100101111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100101111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100110000000000000) && ({row_reg, col_reg}<19'b0100110000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000010010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110000010010101) && ({row_reg, col_reg}<19'b0100110000011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000011000100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100110000011000101)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0100110000011000110)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}==19'b0100110000011000111)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0100110000011001000)) color_data = 12'b000100010100;
		if(({row_reg, col_reg}==19'b0100110000011001001)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==19'b0100110000011001010)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0100110000011001011)) color_data = 12'b000100010011;
		if(({row_reg, col_reg}>=19'b0100110000011001100) && ({row_reg, col_reg}<19'b0100110000011001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100110000011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0100110000011001111) && ({row_reg, col_reg}<19'b0100110000011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100110000011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110000011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100110000011110011) && ({row_reg, col_reg}<19'b0100110000011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000011110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110000011110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100110000011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110000011111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100110000011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110000011111100) && ({row_reg, col_reg}<19'b0100110000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110000011111111) && ({row_reg, col_reg}<19'b0100110000100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110000100000010) && ({row_reg, col_reg}<19'b0100110000100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000100000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110000100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110000100000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0100110000100000111) && ({row_reg, col_reg}<19'b0100110000100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100110000100001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110000100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110000100001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0100110000100001110) && ({row_reg, col_reg}<19'b0100110000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110000100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110000100011001) && ({row_reg, col_reg}<19'b0100110000100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100110000100011100) && ({row_reg, col_reg}<19'b0100110000100011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100110000100011110) && ({row_reg, col_reg}<19'b0100110001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100110001001010001) && ({row_reg, col_reg}<19'b0100110001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100110001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100110001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100110010000000000) && ({row_reg, col_reg}<19'b0100110010011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110010011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0100110010011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100110010011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110010011000100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0100110010011000101)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==19'b0100110010011000110)) color_data = 12'b001000100110;
		if(({row_reg, col_reg}>=19'b0100110010011000111) && ({row_reg, col_reg}<19'b0100110010011001001)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==19'b0100110010011001001)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0100110010011001010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0100110010011001011) && ({row_reg, col_reg}<19'b0100110010011001101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100110010011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110010011001110) && ({row_reg, col_reg}<19'b0100110010011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110010011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100110010011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110010011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100110010011110011) && ({row_reg, col_reg}<19'b0100110010011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110010011110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110010011110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100110010011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110010011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100110010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110010011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110010011111100) && ({row_reg, col_reg}<19'b0100110010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110010011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110010011111111) && ({row_reg, col_reg}<19'b0100110010100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110010100000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110010100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110010100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0100110010100000111) && ({row_reg, col_reg}<19'b0100110010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110010100001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110010100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110010100001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0100110010100001110) && ({row_reg, col_reg}<19'b0100110010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110010100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100110010100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110010100011010) && ({row_reg, col_reg}<19'b0100110011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100110011001010001) && ({row_reg, col_reg}<19'b0100110011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100110011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100110011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100110100000000000) && ({row_reg, col_reg}<19'b0100110100011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110100011000001)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0100110100011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100110100011000011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100110100011000100)) color_data = 12'b000100010100;
		if(({row_reg, col_reg}==19'b0100110100011000101)) color_data = 12'b010000110111;
		if(({row_reg, col_reg}==19'b0100110100011000110)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}==19'b0100110100011000111)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==19'b0100110100011001000)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==19'b0100110100011001001)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0100110100011001010)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0100110100011001011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0100110100011001100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100110100011001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110100011001110)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0100110100011001111) && ({row_reg, col_reg}<19'b0100110100011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110100011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100110100011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110100011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100110100011110011) && ({row_reg, col_reg}<19'b0100110100011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110100011110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110100011110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110100011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110100011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100110100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110100011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110100011111100) && ({row_reg, col_reg}<19'b0100110100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110100011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110100011111111) && ({row_reg, col_reg}<19'b0100110100100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110100100000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110100100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110100100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0100110100100000111) && ({row_reg, col_reg}<19'b0100110100100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110100100001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110100100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110100100001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110100100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110100100001111) && ({row_reg, col_reg}<19'b0100110100100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110100100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100110100100011001) && ({row_reg, col_reg}<19'b0100110101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100110101001010001) && ({row_reg, col_reg}<19'b0100110101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100110101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100110101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100110110000000000) && ({row_reg, col_reg}<19'b0100110110010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110110010010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110110010010101) && ({row_reg, col_reg}<19'b0100110110010010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100110110010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110110010011000) && ({row_reg, col_reg}<19'b0100110110011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110110011000001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0100110110011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100110110011000011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0100110110011000100)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==19'b0100110110011000101)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}==19'b0100110110011000110)) color_data = 12'b011001011011;
		if(({row_reg, col_reg}==19'b0100110110011000111)) color_data = 12'b010101001011;
		if(({row_reg, col_reg}==19'b0100110110011001000)) color_data = 12'b001100011000;
		if(({row_reg, col_reg}==19'b0100110110011001001)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==19'b0100110110011001010)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0100110110011001011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0100110110011001100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100110110011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110110011001110) && ({row_reg, col_reg}<19'b0100110110011010000)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}>=19'b0100110110011010000) && ({row_reg, col_reg}<19'b0100110110011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110110011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100110110011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110110011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100110110011110011) && ({row_reg, col_reg}<19'b0100110110011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110110011110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100110110011110111) && ({row_reg, col_reg}<19'b0100110110011111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110110011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100110110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110110011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110110011111100) && ({row_reg, col_reg}<19'b0100110110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110110011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110110011111111) && ({row_reg, col_reg}<19'b0100110110100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110110100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100110110100000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100110110100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110110100000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0100110110100000111) && ({row_reg, col_reg}<19'b0100110110100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100110110100001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110110100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110110100001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110110100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100110110100001111) && ({row_reg, col_reg}<19'b0100110110100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100110110100011100) && ({row_reg, col_reg}<19'b0100110110100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100110110100100000) && ({row_reg, col_reg}<19'b0100110111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100110111001010001) && ({row_reg, col_reg}<19'b0100110111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100110111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100110111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100111000000000000) && ({row_reg, col_reg}<19'b0100111000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111000010010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100111000010010101) && ({row_reg, col_reg}<19'b0100111000010010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111000010010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100111000010011000) && ({row_reg, col_reg}<19'b0100111000011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111000011000001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0100111000011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111000011000011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100111000011000100)) color_data = 12'b000100010100;
		if(({row_reg, col_reg}==19'b0100111000011000101)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}>=19'b0100111000011000110) && ({row_reg, col_reg}<19'b0100111000011001000)) color_data = 12'b011001011100;
		if(({row_reg, col_reg}==19'b0100111000011001000)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==19'b0100111000011001001)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==19'b0100111000011001010)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0100111000011001011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0100111000011001100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100111000011001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100111000011001110) && ({row_reg, col_reg}<19'b0100111000011010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0100111000011010000) && ({row_reg, col_reg}<19'b0100111000011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111000011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111000011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111000011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100111000011110011) && ({row_reg, col_reg}<19'b0100111000011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111000011110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100111000011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111000011111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100111000011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100111000011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111000011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111000011111100) && ({row_reg, col_reg}<19'b0100111000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111000011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111000011111111) && ({row_reg, col_reg}<19'b0100111000100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111000100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100111000100000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111000100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111000100000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100111000100000111) && ({row_reg, col_reg}<19'b0100111000100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111000100001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100111000100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111000100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100111000100001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100111000100001111) && ({row_reg, col_reg}<19'b0100111000100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100111000100011011) && ({row_reg, col_reg}<19'b0100111000100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111000100011101) && ({row_reg, col_reg}<19'b0100111000111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111000111001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111000111010000) && ({row_reg, col_reg}<19'b0100111001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100111001001010001) && ({row_reg, col_reg}<19'b0100111001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100111001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100111001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100111010000000000) && ({row_reg, col_reg}<19'b0100111010010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010010010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100111010010010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111010010010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100111010010010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100111010010011000) && ({row_reg, col_reg}<19'b0100111010011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010011000011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100111010011000100)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==19'b0100111010011000101)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}==19'b0100111010011000110)) color_data = 12'b011001011100;
		if(({row_reg, col_reg}==19'b0100111010011000111)) color_data = 12'b011001011101;
		if(({row_reg, col_reg}==19'b0100111010011001000)) color_data = 12'b001100101010;
		if(({row_reg, col_reg}==19'b0100111010011001001)) color_data = 12'b001000011000;
		if(({row_reg, col_reg}==19'b0100111010011001010)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==19'b0100111010011001011)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0100111010011001100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0100111010011001101) && ({row_reg, col_reg}<19'b0100111010011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111010011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111010011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100111010011110011) && ({row_reg, col_reg}<19'b0100111010011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010011110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100111010011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111010011111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111010011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111010011111100) && ({row_reg, col_reg}<19'b0100111010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111010011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111010100000001) && ({row_reg, col_reg}<19'b0100111010100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010100000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100111010100000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100111010100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111010100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010100000111) && ({row_reg, col_reg}<19'b0100111010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010100001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100111010100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111010100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100111010100001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100111010100001111) && ({row_reg, col_reg}<19'b0100111010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111010100011011) && ({row_reg, col_reg}<19'b0100111010111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010111000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111010111000011) && ({row_reg, col_reg}<19'b0100111010111001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100111010111001001) && ({row_reg, col_reg}<19'b0100111010111001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100111010111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111010111001100) && ({row_reg, col_reg}<19'b0100111010111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111010111001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111010111010000) && ({row_reg, col_reg}<19'b0100111011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100111011001010001) && ({row_reg, col_reg}<19'b0100111011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100111011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100111011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100111100000000000) && ({row_reg, col_reg}<19'b0100111100010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100010010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111100010010010) && ({row_reg, col_reg}<19'b0100111100010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100010010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100111100010010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111100010010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111100010010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0100111100010011000) && ({row_reg, col_reg}<19'b0100111100011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100111100011000001) && ({row_reg, col_reg}<19'b0100111100011000011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0100111100011000011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100111100011000100)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==19'b0100111100011000101)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}>=19'b0100111100011000110) && ({row_reg, col_reg}<19'b0100111100011001000)) color_data = 12'b011101011101;
		if(({row_reg, col_reg}==19'b0100111100011001000)) color_data = 12'b011001001101;
		if(({row_reg, col_reg}==19'b0100111100011001001)) color_data = 12'b010000111011;
		if(({row_reg, col_reg}==19'b0100111100011001010)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==19'b0100111100011001011)) color_data = 12'b001000100110;
		if(({row_reg, col_reg}==19'b0100111100011001100)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==19'b0100111100011001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100111100011001110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0100111100011001111) && ({row_reg, col_reg}<19'b0100111100011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111100011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111100011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100111100011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100011110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111100011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100011110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111100011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111100011111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111100011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111100011111100) && ({row_reg, col_reg}<19'b0100111100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111100011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111100100000001) && ({row_reg, col_reg}<19'b0100111100100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100100000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100111100100000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111100100000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111100100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100100000111) && ({row_reg, col_reg}<19'b0100111100100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111100100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100100001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100111100100001100) && ({row_reg, col_reg}<19'b0100111100100001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111100100001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100111100100001111) && ({row_reg, col_reg}<19'b0100111100100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111100100011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100111100100100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100111100100100001) && ({row_reg, col_reg}<19'b0100111100100100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100111100100100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0100111100100100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100111100100100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0100111100100100111) && ({row_reg, col_reg}<19'b0100111100111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100111000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0100111100111000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100111100111000100) && ({row_reg, col_reg}<19'b0100111100111001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100111001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111100111001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100111001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0100111100111001100) && ({row_reg, col_reg}<19'b0100111100111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111100111001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111100111010000) && ({row_reg, col_reg}<19'b0100111101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100111101001010001) && ({row_reg, col_reg}<19'b0100111101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100111101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100111101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0100111110000000000) && ({row_reg, col_reg}<19'b0100111110010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110010010001)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0100111110010010010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0100111110010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110010010100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==19'b0100111110010010101)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0100111110010010110)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==19'b0100111110010010111)) color_data = 12'b101110111001;
		if(({row_reg, col_reg}>=19'b0100111110010011000) && ({row_reg, col_reg}<19'b0100111110010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100111110010011101) && ({row_reg, col_reg}<19'b0100111110010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0100111110010100000) && ({row_reg, col_reg}<19'b0100111110011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110011000000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0100111110011000001)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0100111110011000010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0100111110011000011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0100111110011000100)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==19'b0100111110011000101)) color_data = 12'b010001001010;
		if(({row_reg, col_reg}==19'b0100111110011000110)) color_data = 12'b011101101110;
		if(({row_reg, col_reg}==19'b0100111110011000111)) color_data = 12'b011001101110;
		if(({row_reg, col_reg}==19'b0100111110011001000)) color_data = 12'b100001111111;
		if(({row_reg, col_reg}==19'b0100111110011001001)) color_data = 12'b011101111110;
		if(({row_reg, col_reg}==19'b0100111110011001010)) color_data = 12'b011001101100;
		if(({row_reg, col_reg}==19'b0100111110011001011)) color_data = 12'b010101011010;
		if(({row_reg, col_reg}==19'b0100111110011001100)) color_data = 12'b010101011000;
		if(({row_reg, col_reg}==19'b0100111110011001101)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==19'b0100111110011001110)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0100111110011001111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0100111110011010000) && ({row_reg, col_reg}<19'b0100111110011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111110011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111110011110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100111110011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110011110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111110011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110011110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111110011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111110011111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100111110011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111110011111100) && ({row_reg, col_reg}<19'b0100111110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111110011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0100111110100000001) && ({row_reg, col_reg}<19'b0100111110100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110100000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0100111110100000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111110100000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111110100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110100000111) && ({row_reg, col_reg}<19'b0100111110100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0100111110100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110100001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0100111110100001100) && ({row_reg, col_reg}<19'b0100111110100001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111110100001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0100111110100001111) && ({row_reg, col_reg}<19'b0100111110100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110100011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0100111110100011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111110100011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0100111110100100000) && ({row_reg, col_reg}<19'b0100111110100100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111110100100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111110100100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100111110100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111110100101000) && ({row_reg, col_reg}<19'b0100111110111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110111000010)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==19'b0100111110111000011)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==19'b0100111110111000100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=19'b0100111110111000101) && ({row_reg, col_reg}<19'b0100111110111000111)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0100111110111000111)) color_data = 12'b101110111100;
		if(({row_reg, col_reg}>=19'b0100111110111001000) && ({row_reg, col_reg}<19'b0100111110111001010)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0100111110111001010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==19'b0100111110111001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0100111110111001100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0100111110111001101) && ({row_reg, col_reg}<19'b0100111110111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0100111110111001111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0100111110111010000) && ({row_reg, col_reg}<19'b0100111111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0100111111001010001) && ({row_reg, col_reg}<19'b0100111111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0100111111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0100111111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101000000000000000) && ({row_reg, col_reg}<19'b0101000000010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000010010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=19'b0101000000010010001) && ({row_reg, col_reg}<19'b0101000000010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000010010011)) color_data = 12'b010101100010;
		if(({row_reg, col_reg}==19'b0101000000010010100)) color_data = 12'b110111011000;
		if(({row_reg, col_reg}==19'b0101000000010010101)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}>=19'b0101000000010010110) && ({row_reg, col_reg}<19'b0101000000010011000)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}>=19'b0101000000010011000) && ({row_reg, col_reg}<19'b0101000000010011010)) color_data = 12'b001000110000;
		if(({row_reg, col_reg}==19'b0101000000010011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0101000000010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0101000000010011100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101000000010011101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101000000010011110)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101000000010011111)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0101000000010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101000000010100001) && ({row_reg, col_reg}<19'b0101000000011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000011000000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0101000000011000001)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0101000000011000010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101000000011000011)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0101000000011000100)) color_data = 12'b000100101000;
		if(({row_reg, col_reg}==19'b0101000000011000101)) color_data = 12'b001101001100;
		if(({row_reg, col_reg}>=19'b0101000000011000110) && ({row_reg, col_reg}<19'b0101000000011001000)) color_data = 12'b010001011110;
		if(({row_reg, col_reg}==19'b0101000000011001000)) color_data = 12'b010001001110;
		if(({row_reg, col_reg}==19'b0101000000011001001)) color_data = 12'b011001101111;
		if(({row_reg, col_reg}==19'b0101000000011001010)) color_data = 12'b011001111111;
		if(({row_reg, col_reg}==19'b0101000000011001011)) color_data = 12'b010101101100;
		if(({row_reg, col_reg}==19'b0101000000011001100)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==19'b0101000000011001101)) color_data = 12'b010001100111;
		if(({row_reg, col_reg}==19'b0101000000011001110)) color_data = 12'b000100110011;
		if(({row_reg, col_reg}>=19'b0101000000011001111) && ({row_reg, col_reg}<19'b0101000000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000000011110000) && ({row_reg, col_reg}<19'b0101000000011110010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101000000011110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101000000011110011) && ({row_reg, col_reg}<19'b0101000000011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000000011110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101000000011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000000011111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101000000011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101000000011111010) && ({row_reg, col_reg}<19'b0101000000011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000011111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101000000011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000000011111110) && ({row_reg, col_reg}<19'b0101000000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000000100000001) && ({row_reg, col_reg}<19'b0101000000100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000100000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101000000100000100) && ({row_reg, col_reg}<19'b0101000000100000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000000100000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101000000100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101000000100001000) && ({row_reg, col_reg}<19'b0101000000100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101000000100001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101000000100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000000100001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101000000100001111) && ({row_reg, col_reg}<19'b0101000000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000000100010001) && ({row_reg, col_reg}<19'b0101000000100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000000100010011) && ({row_reg, col_reg}<19'b0101000000100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000100011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101000000100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000000100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101000000100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000000100011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000000100011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101000000100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000000100100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101000000100100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101000000100100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101000000100100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0101000000100100101) && ({row_reg, col_reg}<19'b0101000000100100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000000100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000000100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101000000100101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101000000100101010) && ({row_reg, col_reg}<19'b0101000000100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000000100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000000100110000) && ({row_reg, col_reg}<19'b0101000000101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000000101000000) && ({row_reg, col_reg}<19'b0101000000101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000000101000100) && ({row_reg, col_reg}<19'b0101000000101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000000101011001) && ({row_reg, col_reg}<19'b0101000000101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000000101011101) && ({row_reg, col_reg}<19'b0101000000110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000000110111100) && ({row_reg, col_reg}<19'b0101000000110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000000110111110) && ({row_reg, col_reg}<19'b0101000000111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000000111000000) && ({row_reg, col_reg}<19'b0101000000111000010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0101000000111000010)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0101000000111000011)) color_data = 12'b100101111010;
		if(({row_reg, col_reg}==19'b0101000000111000100)) color_data = 12'b110010011100;
		if(({row_reg, col_reg}==19'b0101000000111000101)) color_data = 12'b011101000111;
		if(({row_reg, col_reg}==19'b0101000000111000110)) color_data = 12'b001100000011;
		if(({row_reg, col_reg}==19'b0101000000111000111)) color_data = 12'b010000010100;
		if(({row_reg, col_reg}==19'b0101000000111001000)) color_data = 12'b001100000011;
		if(({row_reg, col_reg}>=19'b0101000000111001001) && ({row_reg, col_reg}<19'b0101000000111001011)) color_data = 12'b111011001111;
		if(({row_reg, col_reg}==19'b0101000000111001011)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==19'b0101000000111001100)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101000000111001101)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0101000000111001110) && ({row_reg, col_reg}<19'b0101000000111010000)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0101000000111010000) && ({row_reg, col_reg}<19'b0101000001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000001001010001) && ({row_reg, col_reg}<19'b0101000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101000001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101000001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101000010000000000) && ({row_reg, col_reg}<19'b0101000010010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010010010000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0101000010010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010010010010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0101000010010010011)) color_data = 12'b100110100100;
		if(({row_reg, col_reg}==19'b0101000010010010100)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}==19'b0101000010010010101)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==19'b0101000010010010110)) color_data = 12'b111111110111;
		if(({row_reg, col_reg}==19'b0101000010010010111)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==19'b0101000010010011000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==19'b0101000010010011001)) color_data = 12'b001101000000;
		if(({row_reg, col_reg}==19'b0101000010010011010)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0101000010010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010010011100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101000010010011101)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101000010010011110)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==19'b0101000010010011111)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==19'b0101000010010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101000010010100001) && ({row_reg, col_reg}<19'b0101000010011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000010011000000) && ({row_reg, col_reg}<19'b0101000010011000010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0101000010011000010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101000010011000011)) color_data = 12'b000000010101;
		if(({row_reg, col_reg}==19'b0101000010011000100)) color_data = 12'b001000111001;
		if(({row_reg, col_reg}==19'b0101000010011000101)) color_data = 12'b010001011101;
		if(({row_reg, col_reg}>=19'b0101000010011000110) && ({row_reg, col_reg}<19'b0101000010011001000)) color_data = 12'b010001011111;
		if(({row_reg, col_reg}==19'b0101000010011001000)) color_data = 12'b010001001111;
		if(({row_reg, col_reg}==19'b0101000010011001001)) color_data = 12'b010101101111;
		if(({row_reg, col_reg}==19'b0101000010011001010)) color_data = 12'b010101111110;
		if(({row_reg, col_reg}==19'b0101000010011001011)) color_data = 12'b001101011011;
		if(({row_reg, col_reg}==19'b0101000010011001100)) color_data = 12'b001001001000;
		if(({row_reg, col_reg}==19'b0101000010011001101)) color_data = 12'b001001000110;
		if(({row_reg, col_reg}==19'b0101000010011001110)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}>=19'b0101000010011001111) && ({row_reg, col_reg}<19'b0101000010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010011110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101000010011110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000010011110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101000010011110011) && ({row_reg, col_reg}<19'b0101000010011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010011110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101000010011110111) && ({row_reg, col_reg}<19'b0101000010011111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000010011111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101000010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000010011111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101000010011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000010100000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101000010100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000010100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010100000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101000010100000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000010100000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000010100000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101000010100000111) && ({row_reg, col_reg}<19'b0101000010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101000010100001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101000010100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000010100001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101000010100001111) && ({row_reg, col_reg}<19'b0101000010100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000010100010011) && ({row_reg, col_reg}<19'b0101000010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101000010100011001) && ({row_reg, col_reg}<19'b0101000010100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000010100011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101000010100011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101000010100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000010100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000010100100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101000010100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000010100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010100100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101000010100100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101000010100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000010100100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101000010100100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101000010100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000010100101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101000010100101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000010100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101000010100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000010100101101) && ({row_reg, col_reg}<19'b0101000010100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101000010100110000) && ({row_reg, col_reg}<19'b0101000010100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000010100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101000010100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000010100111100) && ({row_reg, col_reg}<19'b0101000010101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000010101000110) && ({row_reg, col_reg}<19'b0101000010101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000010101001000) && ({row_reg, col_reg}<19'b0101000010101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000010101011000) && ({row_reg, col_reg}<19'b0101000010101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000010101011111) && ({row_reg, col_reg}<19'b0101000010101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000010101100010) && ({row_reg, col_reg}<19'b0101000010110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000010110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000010110111110) && ({row_reg, col_reg}<19'b0101000010111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000010111000000) && ({row_reg, col_reg}<19'b0101000010111000010)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101000010111000010)) color_data = 12'b010100010101;
		if(({row_reg, col_reg}==19'b0101000010111000011)) color_data = 12'b101110001100;
		if(({row_reg, col_reg}==19'b0101000010111000100)) color_data = 12'b110010001100;
		if(({row_reg, col_reg}==19'b0101000010111000101)) color_data = 12'b011000110110;
		if(({row_reg, col_reg}==19'b0101000010111000110)) color_data = 12'b001100000011;
		if(({row_reg, col_reg}==19'b0101000010111000111)) color_data = 12'b001100000100;
		if(({row_reg, col_reg}==19'b0101000010111001000)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}>=19'b0101000010111001001) && ({row_reg, col_reg}<19'b0101000010111001011)) color_data = 12'b110110101110;
		if(({row_reg, col_reg}==19'b0101000010111001011)) color_data = 12'b010000010100;
		if(({row_reg, col_reg}==19'b0101000010111001100)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101000010111001101)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}>=19'b0101000010111001110) && ({row_reg, col_reg}<19'b0101000010111010000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0101000010111010000) && ({row_reg, col_reg}<19'b0101000011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000011001010001) && ({row_reg, col_reg}<19'b0101000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101000011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101000011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101000100000000000) && ({row_reg, col_reg}<19'b0101000100010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100010010001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0101000100010010010)) color_data = 12'b011101110100;
		if(({row_reg, col_reg}==19'b0101000100010010011)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0101000100010010100)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==19'b0101000100010010101)) color_data = 12'b111011111000;
		if(({row_reg, col_reg}==19'b0101000100010010110)) color_data = 12'b111011110111;
		if(({row_reg, col_reg}==19'b0101000100010010111)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==19'b0101000100010011000)) color_data = 12'b101111010101;
		if(({row_reg, col_reg}==19'b0101000100010011001)) color_data = 12'b100010010011;
		if(({row_reg, col_reg}==19'b0101000100010011010)) color_data = 12'b001100110000;
		if(({row_reg, col_reg}==19'b0101000100010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100010011100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101000100010011101)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0101000100010011110)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==19'b0101000100010011111)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0101000100010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101000100010100001) && ({row_reg, col_reg}<19'b0101000100011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100011000001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0101000100011000010)) color_data = 12'b000000100011;
		if(({row_reg, col_reg}==19'b0101000100011000011)) color_data = 12'b001001000111;
		if(({row_reg, col_reg}==19'b0101000100011000100)) color_data = 12'b010001101100;
		if(({row_reg, col_reg}==19'b0101000100011000101)) color_data = 12'b010101111110;
		if(({row_reg, col_reg}==19'b0101000100011000110)) color_data = 12'b010101101111;
		if(({row_reg, col_reg}==19'b0101000100011000111)) color_data = 12'b010001011111;
		if(({row_reg, col_reg}==19'b0101000100011001000)) color_data = 12'b010001011110;
		if(({row_reg, col_reg}==19'b0101000100011001001)) color_data = 12'b010101101111;
		if(({row_reg, col_reg}==19'b0101000100011001010)) color_data = 12'b010101101101;
		if(({row_reg, col_reg}==19'b0101000100011001011)) color_data = 12'b001001001001;
		if(({row_reg, col_reg}==19'b0101000100011001100)) color_data = 12'b000000100110;
		if(({row_reg, col_reg}==19'b0101000100011001101)) color_data = 12'b000000100100;
		if(({row_reg, col_reg}==19'b0101000100011001110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0101000100011001111) && ({row_reg, col_reg}<19'b0101000100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000100011110000) && ({row_reg, col_reg}<19'b0101000100011110010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000100011110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000100011110011) && ({row_reg, col_reg}<19'b0101000100011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100011110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101000100011110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101000100011111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000100011111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101000100011111010) && ({row_reg, col_reg}<19'b0101000100011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000100100000000) && ({row_reg, col_reg}<19'b0101000100100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100100000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101000100100000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000100100000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000100100000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101000100100000111) && ({row_reg, col_reg}<19'b0101000100100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000100100001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101000100100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000100100001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101000100100001111) && ({row_reg, col_reg}<19'b0101000100100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000100100010011) && ({row_reg, col_reg}<19'b0101000100100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000100100010110) && ({row_reg, col_reg}<19'b0101000100100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000100100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100100011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101000100100011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000100100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000100100011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101000100100011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101000100100011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101000100100100000) && ({row_reg, col_reg}<19'b0101000100100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101000100100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000100100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101000100100101001) && ({row_reg, col_reg}<19'b0101000100100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000100100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101000100100101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101000100100101101) && ({row_reg, col_reg}<19'b0101000100100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101000100100110000) && ({row_reg, col_reg}<19'b0101000100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000100100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101000100100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000100100111100) && ({row_reg, col_reg}<19'b0101000100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000100100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000100101000000) && ({row_reg, col_reg}<19'b0101000100101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000100101011110) && ({row_reg, col_reg}<19'b0101000100101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000100101100010) && ({row_reg, col_reg}<19'b0101000100110111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000100110111111) && ({row_reg, col_reg}<19'b0101000100111000001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0101000100111000001)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0101000100111000010)) color_data = 12'b011101001000;
		if(({row_reg, col_reg}==19'b0101000100111000011)) color_data = 12'b110010001100;
		if(({row_reg, col_reg}==19'b0101000100111000100)) color_data = 12'b101001111010;
		if(({row_reg, col_reg}==19'b0101000100111000101)) color_data = 12'b001100000100;
		if(({row_reg, col_reg}==19'b0101000100111000110)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101000100111000111)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0101000100111001000)) color_data = 12'b001100000100;
		if(({row_reg, col_reg}==19'b0101000100111001001)) color_data = 12'b110010011101;
		if(({row_reg, col_reg}==19'b0101000100111001010)) color_data = 12'b101110001100;
		if(({row_reg, col_reg}==19'b0101000100111001011)) color_data = 12'b001100000011;
		if(({row_reg, col_reg}==19'b0101000100111001100)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101000100111001101)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0101000100111001110)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101000100111001111)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0101000100111010000) && ({row_reg, col_reg}<19'b0101000101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000101001010001) && ({row_reg, col_reg}<19'b0101000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101000101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101000101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101000110000000000) && ({row_reg, col_reg}<19'b0101000110010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110010010000)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==19'b0101000110010010001)) color_data = 12'b011110000101;
		if(({row_reg, col_reg}==19'b0101000110010010010)) color_data = 12'b110011011010;
		if(({row_reg, col_reg}==19'b0101000110010010011)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0101000110010010100)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}==19'b0101000110010010101)) color_data = 12'b110011010110;
		if(({row_reg, col_reg}==19'b0101000110010010110)) color_data = 12'b110011100110;
		if(({row_reg, col_reg}==19'b0101000110010010111)) color_data = 12'b111011111000;
		if(({row_reg, col_reg}==19'b0101000110010011000)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==19'b0101000110010011001)) color_data = 12'b110011010111;
		if(({row_reg, col_reg}==19'b0101000110010011010)) color_data = 12'b010101010010;
		if(({row_reg, col_reg}==19'b0101000110010011011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0101000110010011100)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101000110010011101)) color_data = 12'b000100010100;
		if(({row_reg, col_reg}==19'b0101000110010011110)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==19'b0101000110010011111)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101000110010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101000110010100001) && ({row_reg, col_reg}<19'b0101000110011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110011000001)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}==19'b0101000110011000010)) color_data = 12'b001001000110;
		if(({row_reg, col_reg}==19'b0101000110011000011)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==19'b0101000110011000100)) color_data = 12'b011010001101;
		if(({row_reg, col_reg}==19'b0101000110011000101)) color_data = 12'b011001111110;
		if(({row_reg, col_reg}==19'b0101000110011000110)) color_data = 12'b010101101110;
		if(({row_reg, col_reg}==19'b0101000110011000111)) color_data = 12'b010001001101;
		if(({row_reg, col_reg}==19'b0101000110011001000)) color_data = 12'b010001011110;
		if(({row_reg, col_reg}==19'b0101000110011001001)) color_data = 12'b010101101111;
		if(({row_reg, col_reg}==19'b0101000110011001010)) color_data = 12'b010001101101;
		if(({row_reg, col_reg}==19'b0101000110011001011)) color_data = 12'b000100111000;
		if(({row_reg, col_reg}==19'b0101000110011001100)) color_data = 12'b000000010100;
		if(({row_reg, col_reg}==19'b0101000110011001101)) color_data = 12'b000000010011;
		if(({row_reg, col_reg}==19'b0101000110011001110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0101000110011001111) && ({row_reg, col_reg}<19'b0101000110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000110011110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000110011110011) && ({row_reg, col_reg}<19'b0101000110011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110011110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101000110011110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000110011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000110011111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000110011111010) && ({row_reg, col_reg}<19'b0101000110011111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101000110011111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101000110011111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101000110011111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101000110011111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101000110100000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101000110100000001) && ({row_reg, col_reg}<19'b0101000110100000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101000110100000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101000110100000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000110100000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101000110100000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101000110100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101000110100001000) && ({row_reg, col_reg}<19'b0101000110100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110100001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000110100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000110100001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101000110100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000110100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101000110100010001) && ({row_reg, col_reg}<19'b0101000110100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000110100010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101000110100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000110100010110) && ({row_reg, col_reg}<19'b0101000110100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110100011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101000110100011010) && ({row_reg, col_reg}<19'b0101000110100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000110100011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101000110100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000110100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110100011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101000110100100000) && ({row_reg, col_reg}<19'b0101000110100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000110100100011) && ({row_reg, col_reg}<19'b0101000110100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000110100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000110100101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101000110100101010) && ({row_reg, col_reg}<19'b0101000110100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000110100101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101000110100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000110100101110) && ({row_reg, col_reg}<19'b0101000110100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000110100111101) && ({row_reg, col_reg}<19'b0101000110101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000110101000000) && ({row_reg, col_reg}<19'b0101000110101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000110101010011) && ({row_reg, col_reg}<19'b0101000110101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000110101011100) && ({row_reg, col_reg}<19'b0101000110101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101000110101011110) && ({row_reg, col_reg}<19'b0101000110110111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101000110110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101000110111000000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0101000110111000001)) color_data = 12'b010100100101;
		if(({row_reg, col_reg}==19'b0101000110111000010)) color_data = 12'b100101101010;
		if(({row_reg, col_reg}==19'b0101000110111000011)) color_data = 12'b101110011100;
		if(({row_reg, col_reg}==19'b0101000110111000100)) color_data = 12'b100001011000;
		if(({row_reg, col_reg}>=19'b0101000110111000101) && ({row_reg, col_reg}<19'b0101000110111000111)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101000110111000111)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0101000110111001000)) color_data = 12'b011000110110;
		if(({row_reg, col_reg}==19'b0101000110111001001)) color_data = 12'b110110101101;
		if(({row_reg, col_reg}==19'b0101000110111001010)) color_data = 12'b101001111011;
		if(({row_reg, col_reg}==19'b0101000110111001011)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0101000110111001100)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101000110111001101)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0101000110111001110) && ({row_reg, col_reg}<19'b0101000110111010000)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0101000110111010000) && ({row_reg, col_reg}<19'b0101000111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101000111001010001) && ({row_reg, col_reg}<19'b0101000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101000111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101000111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101001000000000000) && ({row_reg, col_reg}<19'b0101001000010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000010010000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==19'b0101001000010010001)) color_data = 12'b111011101100;
		if(({row_reg, col_reg}==19'b0101001000010010010)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0101001000010010011)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==19'b0101001000010010100)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=19'b0101001000010010101) && ({row_reg, col_reg}<19'b0101001000010010111)) color_data = 12'b110111100111;
		if(({row_reg, col_reg}>=19'b0101001000010010111) && ({row_reg, col_reg}<19'b0101001000010011001)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}==19'b0101001000010011001)) color_data = 12'b100110100101;
		if(({row_reg, col_reg}==19'b0101001000010011010)) color_data = 12'b001101000001;
		if(({row_reg, col_reg}==19'b0101001000010011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000010011100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101001000010011101)) color_data = 12'b000100010100;
		if(({row_reg, col_reg}==19'b0101001000010011110)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==19'b0101001000010011111)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101001000010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101001000010100001) && ({row_reg, col_reg}<19'b0101001000011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000011000001)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}==19'b0101001000011000010)) color_data = 12'b001001000110;
		if(({row_reg, col_reg}==19'b0101001000011000011)) color_data = 12'b010001101001;
		if(({row_reg, col_reg}==19'b0101001000011000100)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==19'b0101001000011000101)) color_data = 12'b001101001010;
		if(({row_reg, col_reg}==19'b0101001000011000110)) color_data = 12'b001000111010;
		if(({row_reg, col_reg}==19'b0101001000011000111)) color_data = 12'b000100101010;
		if(({row_reg, col_reg}==19'b0101001000011001000)) color_data = 12'b010001011101;
		if(({row_reg, col_reg}==19'b0101001000011001001)) color_data = 12'b011001111110;
		if(({row_reg, col_reg}==19'b0101001000011001010)) color_data = 12'b010101101100;
		if(({row_reg, col_reg}==19'b0101001000011001011)) color_data = 12'b000100110111;
		if(({row_reg, col_reg}==19'b0101001000011001100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101001000011001101)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}==19'b0101001000011001110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0101001000011001111) && ({row_reg, col_reg}<19'b0101001000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000011110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001000011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101001000011110011) && ({row_reg, col_reg}<19'b0101001000011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000011110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001000011110111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101001000011111000) && ({row_reg, col_reg}<19'b0101001000011111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001000011111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001000011111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001000011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0101001000011111101) && ({row_reg, col_reg}<19'b0101001000011111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101001000011111111) && ({row_reg, col_reg}<19'b0101001000100000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001000100000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001000100000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001000100000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101001000100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001000100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001000100001010) && ({row_reg, col_reg}<19'b0101001000100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000100001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101001000100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001000100001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001000100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001000100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001000100010001) && ({row_reg, col_reg}<19'b0101001000100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101001000100010011) && ({row_reg, col_reg}<19'b0101001000100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001000100010101) && ({row_reg, col_reg}<19'b0101001000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000100011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101001000100011001) && ({row_reg, col_reg}<19'b0101001000100011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001000100011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001000100011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101001000100011101) && ({row_reg, col_reg}<19'b0101001000100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000100011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001000100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001000100100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001000100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001000100100100) && ({row_reg, col_reg}<19'b0101001000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001000100101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001000100101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101001000100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001000100101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001000100101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001000100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001000100101111) && ({row_reg, col_reg}<19'b0101001000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001000100110111) && ({row_reg, col_reg}<19'b0101001000100111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101001000100111001) && ({row_reg, col_reg}<19'b0101001000100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000100111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001000100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101001000101000000) && ({row_reg, col_reg}<19'b0101001000101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001000101000111) && ({row_reg, col_reg}<19'b0101001000101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101001000101011000) && ({row_reg, col_reg}<19'b0101001000101011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001000101011010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001000101011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101001000101011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001000101011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101001000101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001000101011111) && ({row_reg, col_reg}<19'b0101001000110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001000110111011) && ({row_reg, col_reg}<19'b0101001000110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001000110111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001000110111111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==19'b0101001000111000000)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==19'b0101001000111000001)) color_data = 12'b100101101001;
		if(({row_reg, col_reg}>=19'b0101001000111000010) && ({row_reg, col_reg}<19'b0101001000111000100)) color_data = 12'b110010011100;
		if(({row_reg, col_reg}==19'b0101001000111000100)) color_data = 12'b011101000111;
		if(({row_reg, col_reg}==19'b0101001000111000101)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0101001000111000110)) color_data = 12'b001100000011;
		if(({row_reg, col_reg}==19'b0101001000111000111)) color_data = 12'b011000110110;
		if(({row_reg, col_reg}==19'b0101001000111001000)) color_data = 12'b100101111010;
		if(({row_reg, col_reg}==19'b0101001000111001001)) color_data = 12'b111011001111;
		if(({row_reg, col_reg}==19'b0101001000111001010)) color_data = 12'b101001111010;
		if(({row_reg, col_reg}==19'b0101001000111001011)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}>=19'b0101001000111001100) && ({row_reg, col_reg}<19'b0101001000111001110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0101001000111001110) && ({row_reg, col_reg}<19'b0101001000111010000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0101001000111010000) && ({row_reg, col_reg}<19'b0101001001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101001001001010001) && ({row_reg, col_reg}<19'b0101001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101001001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101001001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101001010000000000) && ({row_reg, col_reg}<19'b0101001010010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010010010000)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}>=19'b0101001010010010001) && ({row_reg, col_reg}<19'b0101001010010010011)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0101001010010010011)) color_data = 12'b111011101011;
		if(({row_reg, col_reg}==19'b0101001010010010100)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0101001010010010101)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==19'b0101001010010010110)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==19'b0101001010010010111)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}==19'b0101001010010011000)) color_data = 12'b011001100001;
		if(({row_reg, col_reg}==19'b0101001010010011001)) color_data = 12'b001100110000;
		if(({row_reg, col_reg}>=19'b0101001010010011010) && ({row_reg, col_reg}<19'b0101001010010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010010011101)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}==19'b0101001010010011110)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==19'b0101001010010011111)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101001010010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101001010010100001) && ({row_reg, col_reg}<19'b0101001010011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010011000001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0101001010011000010)) color_data = 12'b000000100011;
		if(({row_reg, col_reg}==19'b0101001010011000011)) color_data = 12'b000100100101;
		if(({row_reg, col_reg}==19'b0101001010011000100)) color_data = 12'b000000010101;
		if(({row_reg, col_reg}>=19'b0101001010011000101) && ({row_reg, col_reg}<19'b0101001010011000111)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==19'b0101001010011000111)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==19'b0101001010011001000)) color_data = 12'b001100111010;
		if(({row_reg, col_reg}==19'b0101001010011001001)) color_data = 12'b010101101100;
		if(({row_reg, col_reg}==19'b0101001010011001010)) color_data = 12'b010101101011;
		if(({row_reg, col_reg}==19'b0101001010011001011)) color_data = 12'b000100110111;
		if(({row_reg, col_reg}==19'b0101001010011001100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101001010011001101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0101001010011001110) && ({row_reg, col_reg}<19'b0101001010011010000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0101001010011010000) && ({row_reg, col_reg}<19'b0101001010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010011110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001010011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101001010011110011) && ({row_reg, col_reg}<19'b0101001010011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010011110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001010011111000) && ({row_reg, col_reg}<19'b0101001010011111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001010011111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101001010011111011) && ({row_reg, col_reg}<19'b0101001010011111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001010011111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101001010011111111) && ({row_reg, col_reg}<19'b0101001010100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001010100000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001010100000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001010100000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101001010100000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101001010100000101) && ({row_reg, col_reg}<19'b0101001010100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001010100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001010100001010) && ({row_reg, col_reg}<19'b0101001010100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101001010100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001010100001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001010100001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001010100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001010100010001) && ({row_reg, col_reg}<19'b0101001010100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001010100010100) && ({row_reg, col_reg}<19'b0101001010100010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101001010100011000) && ({row_reg, col_reg}<19'b0101001010100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001010100011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101001010100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001010100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001010100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001010100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101001010100100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001010100100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101001010100100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001010100100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101001010100100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001010100100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001010100100111) && ({row_reg, col_reg}<19'b0101001010100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001010100101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101001010100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001010100101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001010100101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101001010100101111) && ({row_reg, col_reg}<19'b0101001010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001010100110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001010100111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101001010100111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101001010100111010) && ({row_reg, col_reg}<19'b0101001010100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001010100111110) && ({row_reg, col_reg}<19'b0101001010101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010101010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001010101010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101001010101011000) && ({row_reg, col_reg}<19'b0101001010101011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001010101011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101001010101011011) && ({row_reg, col_reg}<19'b0101001010101011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001010101011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001010101011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001010101100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001010101100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001010101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001010101100011) && ({row_reg, col_reg}<19'b0101001010110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001010110111011) && ({row_reg, col_reg}<19'b0101001010110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001010110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001010110111111)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==19'b0101001010111000000)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}==19'b0101001010111000001)) color_data = 12'b110010101101;
		if(({row_reg, col_reg}==19'b0101001010111000010)) color_data = 12'b110110101101;
		if(({row_reg, col_reg}==19'b0101001010111000011)) color_data = 12'b101010001011;
		if(({row_reg, col_reg}==19'b0101001010111000100)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==19'b0101001010111000101)) color_data = 12'b010100100101;
		if(({row_reg, col_reg}==19'b0101001010111000110)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==19'b0101001010111000111)) color_data = 12'b101010001011;
		if(({row_reg, col_reg}==19'b0101001010111001000)) color_data = 12'b101110011100;
		if(({row_reg, col_reg}==19'b0101001010111001001)) color_data = 12'b111011001110;
		if(({row_reg, col_reg}==19'b0101001010111001010)) color_data = 12'b100001101001;
		if(({row_reg, col_reg}==19'b0101001010111001011)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0101001010111001100) && ({row_reg, col_reg}<19'b0101001010111001110)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0101001010111001110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0101001010111001111)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0101001010111010000) && ({row_reg, col_reg}<19'b0101001011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101001011001010001) && ({row_reg, col_reg}<19'b0101001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101001011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101001011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101001100000000000) && ({row_reg, col_reg}<19'b0101001100010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100010010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==19'b0101001100010010001)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}>=19'b0101001100010010010) && ({row_reg, col_reg}<19'b0101001100010010100)) color_data = 12'b011110000101;
		if(({row_reg, col_reg}==19'b0101001100010010100)) color_data = 12'b101111001000;
		if(({row_reg, col_reg}==19'b0101001100010010101)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==19'b0101001100010010110)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0101001100010010111)) color_data = 12'b110011011000;
		if(({row_reg, col_reg}>=19'b0101001100010011000) && ({row_reg, col_reg}<19'b0101001100010011010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101001100010011010) && ({row_reg, col_reg}<19'b0101001100010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100010011101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101001100010011110)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101001100010011111)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101001100010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101001100010100001) && ({row_reg, col_reg}<19'b0101001100011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100011000010)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}==19'b0101001100011000011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101001100011000100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101001100011000101)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0101001100011000110)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}>=19'b0101001100011000111) && ({row_reg, col_reg}<19'b0101001100011001001)) color_data = 12'b000000010111;
		if(({row_reg, col_reg}==19'b0101001100011001001)) color_data = 12'b001101001001;
		if(({row_reg, col_reg}==19'b0101001100011001010)) color_data = 12'b010001011010;
		if(({row_reg, col_reg}==19'b0101001100011001011)) color_data = 12'b000100100110;
		if(({row_reg, col_reg}==19'b0101001100011001100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101001100011001101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101001100011001110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0101001100011001111) && ({row_reg, col_reg}<19'b0101001100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101001100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001100011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101001100011110011) && ({row_reg, col_reg}<19'b0101001100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001100011111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101001100011111010) && ({row_reg, col_reg}<19'b0101001100011111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101001100011111100) && ({row_reg, col_reg}<19'b0101001100011111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101001100011111110) && ({row_reg, col_reg}<19'b0101001100100000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001100100000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001100100000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001100100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001100100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001100100000101) && ({row_reg, col_reg}<19'b0101001100100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001100100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001100100001010) && ({row_reg, col_reg}<19'b0101001100100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001100100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001100100001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001100100001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101001100100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001100100010001) && ({row_reg, col_reg}<19'b0101001100100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001100100010100) && ({row_reg, col_reg}<19'b0101001100100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001100100010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101001100100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001100100011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001100100011010) && ({row_reg, col_reg}<19'b0101001100100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001100100011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001100100011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101001100100100000) && ({row_reg, col_reg}<19'b0101001100100100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001100100100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101001100100100100) && ({row_reg, col_reg}<19'b0101001100100100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001100100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001100100100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001100100101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101001100100101001) && ({row_reg, col_reg}<19'b0101001100100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101001100100101100) && ({row_reg, col_reg}<19'b0101001100100101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001100100101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101001100100101111) && ({row_reg, col_reg}<19'b0101001100100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001100100110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101001100100110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001100100111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001100100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001100100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001100100111100) && ({row_reg, col_reg}<19'b0101001100100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001100100111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101001100101000000) && ({row_reg, col_reg}<19'b0101001100101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001100101000010) && ({row_reg, col_reg}<19'b0101001100101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001100101000100) && ({row_reg, col_reg}<19'b0101001100101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001100101010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001100101010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001100101010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101001100101011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0101001100101011001) && ({row_reg, col_reg}<19'b0101001100101011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101001100101011011) && ({row_reg, col_reg}<19'b0101001100101011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001100101011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001100101100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001100101100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101001100101100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001100101100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001100101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001100101100101) && ({row_reg, col_reg}<19'b0101001100110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001100110111011) && ({row_reg, col_reg}<19'b0101001100110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001100110111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001100110111111)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==19'b0101001100111000000)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0101001100111000001)) color_data = 12'b110010101101;
		if(({row_reg, col_reg}==19'b0101001100111000010)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0101001100111000011)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==19'b0101001100111000100)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0101001100111000101)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}==19'b0101001100111000110)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0101001100111000111)) color_data = 12'b110010111101;
		if(({row_reg, col_reg}==19'b0101001100111001000)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}==19'b0101001100111001001)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0101001100111001010)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==19'b0101001100111001011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0101001100111001100)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==19'b0101001100111001101)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0101001100111001110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0101001100111001111)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=19'b0101001100111010000) && ({row_reg, col_reg}<19'b0101001101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101001101001010001) && ({row_reg, col_reg}<19'b0101001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101001101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101001101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101001110000000000) && ({row_reg, col_reg}<19'b0101001110010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110010010011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0101001110010010100)) color_data = 12'b100110010110;
		if(({row_reg, col_reg}==19'b0101001110010010101)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==19'b0101001110010010110)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==19'b0101001110010010111)) color_data = 12'b100010010101;
		if(({row_reg, col_reg}==19'b0101001110010011000)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0101001110010011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0101001110010011010)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==19'b0101001110010011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001110010011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001110010011101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101001110010011110) && ({row_reg, col_reg}<19'b0101001110010100000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0101001110010100000) && ({row_reg, col_reg}<19'b0101001110011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110011000001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0101001110011000010)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}==19'b0101001110011000011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101001110011000100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101001110011000101)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101001110011000110)) color_data = 12'b000100100110;
		if(({row_reg, col_reg}==19'b0101001110011000111)) color_data = 12'b001101001001;
		if(({row_reg, col_reg}==19'b0101001110011001000)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0101001110011001001)) color_data = 12'b001000110111;
		if(({row_reg, col_reg}==19'b0101001110011001010)) color_data = 12'b010001001000;
		if(({row_reg, col_reg}==19'b0101001110011001011)) color_data = 12'b000100100100;
		if(({row_reg, col_reg}>=19'b0101001110011001100) && ({row_reg, col_reg}<19'b0101001110011001110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101001110011001110) && ({row_reg, col_reg}<19'b0101001110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101001110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101001110011110011) && ({row_reg, col_reg}<19'b0101001110011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001110011110110) && ({row_reg, col_reg}<19'b0101001110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001110011111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001110011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001110011111100) && ({row_reg, col_reg}<19'b0101001110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101001110100000000) && ({row_reg, col_reg}<19'b0101001110100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001110100000010) && ({row_reg, col_reg}<19'b0101001110100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001110100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001110100000110) && ({row_reg, col_reg}<19'b0101001110100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001110100001010) && ({row_reg, col_reg}<19'b0101001110100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001110100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110100001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001110100001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101001110100010000) && ({row_reg, col_reg}<19'b0101001110100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001110100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001110100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001110100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001110100011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101001110100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101001110100011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001110100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001110100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101001110100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110100100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001110100100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110100100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001110100100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101001110100100100) && ({row_reg, col_reg}<19'b0101001110100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110100100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001110100101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101001110100101001) && ({row_reg, col_reg}<19'b0101001110100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001110100101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101001110100101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001110100101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101001110100101111) && ({row_reg, col_reg}<19'b0101001110100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001110100110010) && ({row_reg, col_reg}<19'b0101001110100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101001110100110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101001110100110111) && ({row_reg, col_reg}<19'b0101001110100111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110100111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001110100111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101001110100111100) && ({row_reg, col_reg}<19'b0101001110100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110100111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101001110100111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101001110101000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001110101000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001110101000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101001110101000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001110101000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101001110101000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101001110101000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001110101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001110101001000) && ({row_reg, col_reg}<19'b0101001110101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101001110101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001110101010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001110101010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110101011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101001110101011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001110101011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001110101011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001110101011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001110101011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001110101011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001110101011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101001110101100000) && ({row_reg, col_reg}<19'b0101001110101100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110101100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101001110101100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101001110101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101001110101100101) && ({row_reg, col_reg}<19'b0101001110110111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110110111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101001110110111011) && ({row_reg, col_reg}<19'b0101001110110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101001110110111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101001110110111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101001110111000000)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==19'b0101001110111000001)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==19'b0101001110111000010)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==19'b0101001110111000011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0101001110111000100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101001110111000101)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0101001110111000110)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0101001110111000111)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0101001110111001000)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0101001110111001001)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==19'b0101001110111001010)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==19'b0101001110111001011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101001110111001100)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0101001110111001101)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0101001110111001110)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101001110111001111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0101001110111010000) && ({row_reg, col_reg}<19'b0101001111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101001111001010001) && ({row_reg, col_reg}<19'b0101001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101001111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101001111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101010000000000000) && ({row_reg, col_reg}<19'b0101010000010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000010010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0101010000010010010) && ({row_reg, col_reg}<19'b0101010000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000010010100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==19'b0101010000010010101)) color_data = 12'b110011011010;
		if(({row_reg, col_reg}==19'b0101010000010010110)) color_data = 12'b111011111100;
		if(({row_reg, col_reg}==19'b0101010000010010111)) color_data = 12'b101010111000;
		if(({row_reg, col_reg}>=19'b0101010000010011000) && ({row_reg, col_reg}<19'b0101010000010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010000010011101) && ({row_reg, col_reg}<19'b0101010000010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101010000010100000) && ({row_reg, col_reg}<19'b0101010000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000011000011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101010000011000100) && ({row_reg, col_reg}<19'b0101010000011000110)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0101010000011000110) && ({row_reg, col_reg}<19'b0101010000011001010)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}>=19'b0101010000011001010) && ({row_reg, col_reg}<19'b0101010000011001100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101010000011001100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101010000011001101) && ({row_reg, col_reg}<19'b0101010000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101010000011110011) && ({row_reg, col_reg}<19'b0101010000011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010000011110110) && ({row_reg, col_reg}<19'b0101010000011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010000011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010000011111010) && ({row_reg, col_reg}<19'b0101010000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010000011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010000100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010000100000001) && ({row_reg, col_reg}<19'b0101010000100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010000100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010000100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010000100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101010000100010000) && ({row_reg, col_reg}<19'b0101010000100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000100010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010000100010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010000100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000100011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010000100011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010000100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010000100011011) && ({row_reg, col_reg}<19'b0101010000100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000100011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010000100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000100100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010000100100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101010000100100010) && ({row_reg, col_reg}<19'b0101010000100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000100100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010000100100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010000100100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101010000100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010000100101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010000100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000100101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010000100101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101010000100101111) && ({row_reg, col_reg}<19'b0101010000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000100110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101010000100110011) && ({row_reg, col_reg}<19'b0101010000100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000100110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010000100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000100110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010000100111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010000100111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010000100111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000100111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010000100111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101010000100111110) && ({row_reg, col_reg}<19'b0101010000101000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101010000101000000) && ({row_reg, col_reg}<19'b0101010000101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000101000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010000101000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010000101001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101010000101001001) && ({row_reg, col_reg}<19'b0101010000101001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010000101001101) && ({row_reg, col_reg}<19'b0101010000101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010000101001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101010000101010000) && ({row_reg, col_reg}<19'b0101010000101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010000101010010) && ({row_reg, col_reg}<19'b0101010000101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101010000101010101) && ({row_reg, col_reg}<19'b0101010000101010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000101010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010000101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010000101011010) && ({row_reg, col_reg}<19'b0101010000101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000101011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101010000101011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010000101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000101100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010000101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010000101100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010000101100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000101100100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010000101100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010000101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101010000101101000) && ({row_reg, col_reg}<19'b0101010000101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010000101101011) && ({row_reg, col_reg}<19'b0101010000101101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010000101110000) && ({row_reg, col_reg}<19'b0101010000111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010000111000000)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==19'b0101010000111000001)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0101010000111000010)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0101010000111000011) && ({row_reg, col_reg}<19'b0101010000111000101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0101010000111000101)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0101010000111000110)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0101010000111000111)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=19'b0101010000111001000) && ({row_reg, col_reg}<19'b0101010001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010001001010001) && ({row_reg, col_reg}<19'b0101010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101010001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101010001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101010010000000000) && ({row_reg, col_reg}<19'b0101010010010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010010010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0101010010010010010) && ({row_reg, col_reg}<19'b0101010010010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010010010100)) color_data = 12'b010001010011;
		if(({row_reg, col_reg}==19'b0101010010010010101)) color_data = 12'b110011011011;
		if(({row_reg, col_reg}==19'b0101010010010010110)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0101010010010010111)) color_data = 12'b101111001010;
		if(({row_reg, col_reg}>=19'b0101010010010011000) && ({row_reg, col_reg}<19'b0101010010010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010010010011110) && ({row_reg, col_reg}<19'b0101010010010100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101010010010100000) && ({row_reg, col_reg}<19'b0101010010011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010010011000011) && ({row_reg, col_reg}<19'b0101010010011000110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101010010011000110) && ({row_reg, col_reg}<19'b0101010010011001010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0101010010011001010) && ({row_reg, col_reg}<19'b0101010010011001101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101010010011001101) && ({row_reg, col_reg}<19'b0101010010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101010010011110011) && ({row_reg, col_reg}<19'b0101010010011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010010011110110) && ({row_reg, col_reg}<19'b0101010010100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010010100000101) && ({row_reg, col_reg}<19'b0101010010100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010010100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010010100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101010010100010000) && ({row_reg, col_reg}<19'b0101010010100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010010100010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010010100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010100011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010010100011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010010100011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101010010100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010010100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010010100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010100100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010010100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101010010100100010) && ({row_reg, col_reg}<19'b0101010010100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010010100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010010100100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101010010100100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010010100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010100101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010010100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010010100101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010010100101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010010100101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101010010100101111) && ({row_reg, col_reg}<19'b0101010010100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010010100110011) && ({row_reg, col_reg}<19'b0101010010100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010010100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010100110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010010100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010010100111010) && ({row_reg, col_reg}<19'b0101010010100111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010100111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010010101000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010010101000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101010010101000010) && ({row_reg, col_reg}<19'b0101010010101000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010010101000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010010101000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101010010101000110) && ({row_reg, col_reg}<19'b0101010010101001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010101001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101010010101001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010010101001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101010010101001011) && ({row_reg, col_reg}<19'b0101010010101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010010101010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101010010101010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010010101010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010010101010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010010101010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101010010101011000) && ({row_reg, col_reg}<19'b0101010010101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010010101011101) && ({row_reg, col_reg}<19'b0101010010101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010010101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010101100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010010101100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101010010101100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101010010101100011) && ({row_reg, col_reg}<19'b0101010010101100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010010101100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010010101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101010010101100111) && ({row_reg, col_reg}<19'b0101010010111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010111000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010010111000001)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0101010010111000010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0101010010111000011) && ({row_reg, col_reg}<19'b0101010010111000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010010111000101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0101010010111000110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0101010010111000111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0101010010111001000) && ({row_reg, col_reg}<19'b0101010011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010011001010001) && ({row_reg, col_reg}<19'b0101010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101010011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101010011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101010100000000000) && ({row_reg, col_reg}<19'b0101010100010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100010010001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101010100010010010) && ({row_reg, col_reg}<19'b0101010100010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100010010100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==19'b0101010100010010101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==19'b0101010100010010110)) color_data = 12'b101010111001;
		if(({row_reg, col_reg}==19'b0101010100010010111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=19'b0101010100010011000) && ({row_reg, col_reg}<19'b0101010100011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010100011000101) && ({row_reg, col_reg}<19'b0101010100011001011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101010100011001011) && ({row_reg, col_reg}<19'b0101010100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101010100011110011) && ({row_reg, col_reg}<19'b0101010100011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010100011110110) && ({row_reg, col_reg}<19'b0101010100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010100100000001) && ({row_reg, col_reg}<19'b0101010100100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010100100000100) && ({row_reg, col_reg}<19'b0101010100100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010100100000110) && ({row_reg, col_reg}<19'b0101010100100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010100100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010100100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010100100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101010100100010000) && ({row_reg, col_reg}<19'b0101010100100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100100010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010100100010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100100010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101010100100011000) && ({row_reg, col_reg}<19'b0101010100100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100100011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010100100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101010100100011111) && ({row_reg, col_reg}<19'b0101010100100100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010100100100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101010100100100011) && ({row_reg, col_reg}<19'b0101010100100100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101010100100100111) && ({row_reg, col_reg}<19'b0101010100100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100100101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101010100100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010100100101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010100100101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101010100100101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101010100100101111) && ({row_reg, col_reg}<19'b0101010100100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010100100110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101010100100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100100110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010100100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100100111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010100100111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101010100100111011) && ({row_reg, col_reg}<19'b0101010100100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010100100111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010100101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010100101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010100101000010) && ({row_reg, col_reg}<19'b0101010100101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100101000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010100101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010100101000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010100101000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101010100101001000) && ({row_reg, col_reg}<19'b0101010100101001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100101001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010100101001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101010100101001100) && ({row_reg, col_reg}<19'b0101010100101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100101010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010100101010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010100101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100101010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010100101010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101010100101010111) && ({row_reg, col_reg}<19'b0101010100101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100101100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010100101100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010100101100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010100101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100101100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101010100101100111) && ({row_reg, col_reg}<19'b0101010100111000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100111000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010100111000001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0101010100111000010) && ({row_reg, col_reg}<19'b0101010100111000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010100111000110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0101010100111000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010100111001000) && ({row_reg, col_reg}<19'b0101010101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010101001010001) && ({row_reg, col_reg}<19'b0101010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101010101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101010101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101010110000000000) && ({row_reg, col_reg}<19'b0101010110010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110010010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110010010010) && ({row_reg, col_reg}<19'b0101010110010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010110010010101) && ({row_reg, col_reg}<19'b0101010110010010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010110010010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110010011000) && ({row_reg, col_reg}<19'b0101010110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101010110011110011) && ({row_reg, col_reg}<19'b0101010110011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110011110110) && ({row_reg, col_reg}<19'b0101010110100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010110100000110) && ({row_reg, col_reg}<19'b0101010110100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110100001000) && ({row_reg, col_reg}<19'b0101010110100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010110100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010110100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010110100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101010110100010000) && ({row_reg, col_reg}<19'b0101010110100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010110100010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010110100010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110100010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101010110100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110100011001) && ({row_reg, col_reg}<19'b0101010110100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110100011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101010110100011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010110100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101010110100100000) && ({row_reg, col_reg}<19'b0101010110100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010110100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010110100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110100101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010110100101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010110100101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101010110100101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101010110100101111) && ({row_reg, col_reg}<19'b0101010110100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110100110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010110100110101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010110100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110100110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010110100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110100111001) && ({row_reg, col_reg}<19'b0101010110100111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101010110100111011) && ({row_reg, col_reg}<19'b0101010110100111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010110100111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101010110100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110100111111) && ({row_reg, col_reg}<19'b0101010110101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110101000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110101000110) && ({row_reg, col_reg}<19'b0101010110101001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010110101001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101010110101001001) && ({row_reg, col_reg}<19'b0101010110101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110101001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101010110101001100) && ({row_reg, col_reg}<19'b0101010110101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010110101001110) && ({row_reg, col_reg}<19'b0101010110101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110101010000) && ({row_reg, col_reg}<19'b0101010110101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110101010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101010110101010011) && ({row_reg, col_reg}<19'b0101010110101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101010110101010110) && ({row_reg, col_reg}<19'b0101010110101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101010110101011001) && ({row_reg, col_reg}<19'b0101010110101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110101011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101010110101011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101010110101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101010110101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101010110101100000) && ({row_reg, col_reg}<19'b0101010110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101010110101100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101010110101100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010110101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110101100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101010110101100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101010110101101000) && ({row_reg, col_reg}<19'b0101010111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101010111001010001) && ({row_reg, col_reg}<19'b0101010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101010111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101010111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101011000000000000) && ({row_reg, col_reg}<19'b0101011000010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000010010001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101011000010010010) && ({row_reg, col_reg}<19'b0101011000010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011000010010101) && ({row_reg, col_reg}<19'b0101011000010010111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101011000010010111) && ({row_reg, col_reg}<19'b0101011000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101011000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101011000011110011) && ({row_reg, col_reg}<19'b0101011000011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011000011110110) && ({row_reg, col_reg}<19'b0101011000011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011000011111000) && ({row_reg, col_reg}<19'b0101011000011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011000011111010) && ({row_reg, col_reg}<19'b0101011000011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011000100000000) && ({row_reg, col_reg}<19'b0101011000100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000100000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011000100000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011000100000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101011000100000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011000100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011000100000111) && ({row_reg, col_reg}<19'b0101011000100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011000100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011000100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011000100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101011000100010000) && ({row_reg, col_reg}<19'b0101011000100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000100010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011000100010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011000100010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000100010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101011000100011000) && ({row_reg, col_reg}<19'b0101011000100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000100011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011000100011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101011000100100000) && ({row_reg, col_reg}<19'b0101011000100100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011000100100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101011000100101000) && ({row_reg, col_reg}<19'b0101011000100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011000100101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000100101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011000100101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101011000100101111) && ({row_reg, col_reg}<19'b0101011000100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000100110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011000100110101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011000100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000100110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011000100111000) && ({row_reg, col_reg}<19'b0101011000100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011000100111101) && ({row_reg, col_reg}<19'b0101011000100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011000100111111) && ({row_reg, col_reg}<19'b0101011000101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011000101000011) && ({row_reg, col_reg}<19'b0101011000101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000101001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011000101001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000101001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011000101001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011000101001101) && ({row_reg, col_reg}<19'b0101011000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000101001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011000101010000) && ({row_reg, col_reg}<19'b0101011000101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000101010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011000101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011000101010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101011000101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011000101011000) && ({row_reg, col_reg}<19'b0101011000101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000101011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011000101011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101011000101011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011000101011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101011000101011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011000101011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101011000101100000) && ({row_reg, col_reg}<19'b0101011000101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011000101100010) && ({row_reg, col_reg}<19'b0101011000101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011000101100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011000101100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011000101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000101100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101011000101101000) && ({row_reg, col_reg}<19'b0101011000101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011000101101100) && ({row_reg, col_reg}<19'b0101011000101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011000101101110) && ({row_reg, col_reg}<19'b0101011001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011001001010001) && ({row_reg, col_reg}<19'b0101011001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101011001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101011001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101011010000000000) && ({row_reg, col_reg}<19'b0101011010010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010010010100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101011010010010101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0101011010010010110)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0101011010010010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==19'b0101011010010011000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101011010010011001) && ({row_reg, col_reg}<19'b0101011010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101011010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101011010011110011) && ({row_reg, col_reg}<19'b0101011010011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010011110110) && ({row_reg, col_reg}<19'b0101011010011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011010011111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011010011111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101011010100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011010100000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101011010100000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101011010100000011) && ({row_reg, col_reg}<19'b0101011010100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010100000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011010100000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011010100001000) && ({row_reg, col_reg}<19'b0101011010100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011010100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011010100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011010100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010100010001) && ({row_reg, col_reg}<19'b0101011010100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010100010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101011010100010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011010100010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010100010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101011010100011000) && ({row_reg, col_reg}<19'b0101011010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011010100011010) && ({row_reg, col_reg}<19'b0101011010100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011010100011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010100011101) && ({row_reg, col_reg}<19'b0101011010100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011010100100001) && ({row_reg, col_reg}<19'b0101011010100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010100100011) && ({row_reg, col_reg}<19'b0101011010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011010100100101) && ({row_reg, col_reg}<19'b0101011010100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010100100111) && ({row_reg, col_reg}<19'b0101011010100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010100101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011010100101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011010100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010100101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011010100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010100101111) && ({row_reg, col_reg}<19'b0101011010100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011010100110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011010100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010100110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011010100111000) && ({row_reg, col_reg}<19'b0101011010100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010100111110) && ({row_reg, col_reg}<19'b0101011010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011010101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010101000010) && ({row_reg, col_reg}<19'b0101011010101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010101000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011010101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010101001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101011010101001010) && ({row_reg, col_reg}<19'b0101011010101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010101001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101011010101001101) && ({row_reg, col_reg}<19'b0101011010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011010101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011010101010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011010101010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011010101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011010101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011010101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011010101011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011010101011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101011010101011100) && ({row_reg, col_reg}<19'b0101011010101100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010101100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011010101100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011010101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011010101100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101011010101100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011010101100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010101101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011010101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010101101010) && ({row_reg, col_reg}<19'b0101011010101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011010101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011010101101110) && ({row_reg, col_reg}<19'b0101011011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011011001010001) && ({row_reg, col_reg}<19'b0101011011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101011011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101011011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101011100000000000) && ({row_reg, col_reg}<19'b0101011100010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100010010011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101011100010010100) && ({row_reg, col_reg}<19'b0101011100010010110)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0101011100010010110)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0101011100010010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=19'b0101011100010011000) && ({row_reg, col_reg}<19'b0101011100010011010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101011100010011010) && ({row_reg, col_reg}<19'b0101011100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101011100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101011100011110011) && ({row_reg, col_reg}<19'b0101011100011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011100011110110) && ({row_reg, col_reg}<19'b0101011100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011100011111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011100011111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101011100011111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011100011111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101011100011111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011100100000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101011100100000001) && ({row_reg, col_reg}<19'b0101011100100000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100100000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011100100000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101011100100001000) && ({row_reg, col_reg}<19'b0101011100100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011100100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011100100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011100100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011100100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011100100010001) && ({row_reg, col_reg}<19'b0101011100100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100100010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101011100100010101) && ({row_reg, col_reg}<19'b0101011100100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100100010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101011100100011000) && ({row_reg, col_reg}<19'b0101011100100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011100100011010) && ({row_reg, col_reg}<19'b0101011100100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011100100011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011100100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100100011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011100100011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011100100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011100100100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011100100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011100100100011) && ({row_reg, col_reg}<19'b0101011100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011100100100101) && ({row_reg, col_reg}<19'b0101011100100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011100100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011100100101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011100100101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011100100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100100101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011100100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011100100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011100100110000) && ({row_reg, col_reg}<19'b0101011100100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011100100110011) && ({row_reg, col_reg}<19'b0101011100100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100100110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101011100100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100100110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101011100100111000) && ({row_reg, col_reg}<19'b0101011100100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011100100111010) && ({row_reg, col_reg}<19'b0101011100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011100101000000) && ({row_reg, col_reg}<19'b0101011100101000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011100101000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101011100101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011100101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011100101000110) && ({row_reg, col_reg}<19'b0101011100101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011100101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100101001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011100101001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011100101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100101001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011100101001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011100101001110) && ({row_reg, col_reg}<19'b0101011100101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100101010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101011100101010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011100101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011100101010101) && ({row_reg, col_reg}<19'b0101011100101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011100101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100101011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011100101011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011100101011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101011100101011100) && ({row_reg, col_reg}<19'b0101011100101011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101011100101011110) && ({row_reg, col_reg}<19'b0101011100101100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011100101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011100101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011100101100011) && ({row_reg, col_reg}<19'b0101011100101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100101100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101011100101100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011100101100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100101101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101011100101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011100101101010) && ({row_reg, col_reg}<19'b0101011100101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011100101101101) && ({row_reg, col_reg}<19'b0101011100101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011100101101111) && ({row_reg, col_reg}<19'b0101011100111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011100111000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101011100111000100) && ({row_reg, col_reg}<19'b0101011101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011101001010001) && ({row_reg, col_reg}<19'b0101011101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101011101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101011101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101011110000000000) && ({row_reg, col_reg}<19'b0101011110010010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011110010010011) && ({row_reg, col_reg}<19'b0101011110010011001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101011110010011001) && ({row_reg, col_reg}<19'b0101011110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110011110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101011110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101011110011110011) && ({row_reg, col_reg}<19'b0101011110011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011110011110110) && ({row_reg, col_reg}<19'b0101011110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011110011111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101011110011111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011110011111100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011110011111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101011110011111110) && ({row_reg, col_reg}<19'b0101011110100000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110100000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011110100000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011110100000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011110100000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101011110100000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011110100000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101011110100000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011110100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0101011110100001000) && ({row_reg, col_reg}<19'b0101011110100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011110100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011110100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011110100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011110100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011110100010001) && ({row_reg, col_reg}<19'b0101011110100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110100010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101011110100010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110100010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011110100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011110100011000) && ({row_reg, col_reg}<19'b0101011110100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011110100011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011110100011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011110100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101011110100100001) && ({row_reg, col_reg}<19'b0101011110100100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0101011110100100011) && ({row_reg, col_reg}<19'b0101011110100100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011110100100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011110100100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011110100100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101011110100101000) && ({row_reg, col_reg}<19'b0101011110100101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101011110100101010) && ({row_reg, col_reg}<19'b0101011110100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110100101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011110100101101) && ({row_reg, col_reg}<19'b0101011110100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110100101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101011110100110000) && ({row_reg, col_reg}<19'b0101011110100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110100110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011110100110011) && ({row_reg, col_reg}<19'b0101011110100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110100110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101011110100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110100110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101011110100111000) && ({row_reg, col_reg}<19'b0101011110100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110100111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011110100111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011110100111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011110101000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101011110101000001) && ({row_reg, col_reg}<19'b0101011110101000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110101000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011110101000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011110101000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011110101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110101001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101011110101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110101001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101011110101001011) && ({row_reg, col_reg}<19'b0101011110101001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110101001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101011110101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011110101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110101010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101011110101010010) && ({row_reg, col_reg}<19'b0101011110101010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101011110101010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101011110101010101) && ({row_reg, col_reg}<19'b0101011110101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110101011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101011110101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110101011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101011110101011100) && ({row_reg, col_reg}<19'b0101011110101011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101011110101011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011110101011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101011110101100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110101100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101011110101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101011110101100011) && ({row_reg, col_reg}<19'b0101011110101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101011110101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101011110101100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011110101100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011110101101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101011110101101010) && ({row_reg, col_reg}<19'b0101011110101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011110101101101) && ({row_reg, col_reg}<19'b0101011110101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101011110101101111) && ({row_reg, col_reg}<19'b0101011110111000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011110111000010) && ({row_reg, col_reg}<19'b0101011110111000110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101011110111000110) && ({row_reg, col_reg}<19'b0101011111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101011111001010001) && ({row_reg, col_reg}<19'b0101011111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101011111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101011111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101100000000000000) && ({row_reg, col_reg}<19'b0101100000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000011110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101100000011110011) && ({row_reg, col_reg}<19'b0101100000011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000011111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101100000011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000011111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100000011111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100000011111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101100000011111111) && ({row_reg, col_reg}<19'b0101100000100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100000100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100000100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101100000100000110) && ({row_reg, col_reg}<19'b0101100000100001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000100001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101100000100001001) && ({row_reg, col_reg}<19'b0101100000100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100000100001011) && ({row_reg, col_reg}<19'b0101100000100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100000100001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100000100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101100000100010000) && ({row_reg, col_reg}<19'b0101100000100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100000100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101100000100010101) && ({row_reg, col_reg}<19'b0101100000100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101100000100011010) && ({row_reg, col_reg}<19'b0101100000100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100000100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101100000100011110) && ({row_reg, col_reg}<19'b0101100000100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101100000100100001) && ({row_reg, col_reg}<19'b0101100000100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000100101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100000100101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100000100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100000100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100000100101101) && ({row_reg, col_reg}<19'b0101100000100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100000100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101100000100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000100110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100000100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100000100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100000100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000100111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101100000100111101) && ({row_reg, col_reg}<19'b0101100000100111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000100111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101100000101000000) && ({row_reg, col_reg}<19'b0101100000101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000101000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100000101000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101100000101000100) && ({row_reg, col_reg}<19'b0101100000101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000101000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100000101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000101001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100000101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000101001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100000101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100000101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000101001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100000101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000101001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100000101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000101010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101100000101010100) && ({row_reg, col_reg}<19'b0101100000101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100000101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000101011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101100000101011001) && ({row_reg, col_reg}<19'b0101100000101011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000101011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100000101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100000101011101) && ({row_reg, col_reg}<19'b0101100000101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100000101100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100000101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000101100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100000101100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101100000101100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100000101100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000101101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100000101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101100000101101010) && ({row_reg, col_reg}<19'b0101100000101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100000101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100000101101111) && ({row_reg, col_reg}<19'b0101100000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100000110010100) && ({row_reg, col_reg}<19'b0101100000110010110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0101100000110010110)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0101100000110010111)) color_data = 12'b000100110000;
		if(({row_reg, col_reg}>=19'b0101100000110011000) && ({row_reg, col_reg}<19'b0101100000110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100000110011101) && ({row_reg, col_reg}<19'b0101100000110100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101100000110100000) && ({row_reg, col_reg}<19'b0101100001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100001001010001) && ({row_reg, col_reg}<19'b0101100001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101100001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101100001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101100010000000000) && ({row_reg, col_reg}<19'b0101100010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010011110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101100010011110011) && ({row_reg, col_reg}<19'b0101100010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010011111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100010011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010011111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100010011111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100010011111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101100010011111111) && ({row_reg, col_reg}<19'b0101100010100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101100010100000110) && ({row_reg, col_reg}<19'b0101100010100001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010100001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101100010100001001) && ({row_reg, col_reg}<19'b0101100010100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010100001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100010100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101100010100010000) && ({row_reg, col_reg}<19'b0101100010100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101100010100010101) && ({row_reg, col_reg}<19'b0101100010100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101100010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010100011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100010100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100010100011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101100010100100000) && ({row_reg, col_reg}<19'b0101100010100100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101100010100100011) && ({row_reg, col_reg}<19'b0101100010100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100010100100110) && ({row_reg, col_reg}<19'b0101100010100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100010100101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010100101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100010100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101100010100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100010100101100) && ({row_reg, col_reg}<19'b0101100010100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101100010100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010100110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101100010100111000) && ({row_reg, col_reg}<19'b0101100010100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100010100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010100111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100010100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010101000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101100010101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010101000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010101000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100010101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010101000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100010101000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100010101001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101100010101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010101001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100010101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010101010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100010101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010101010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101100010101010100) && ({row_reg, col_reg}<19'b0101100010101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100010101011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010101011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100010101011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101100010101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100010101011101) && ({row_reg, col_reg}<19'b0101100010101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010101100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100010101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010101100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100010101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010101100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101100010101100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010101101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100010101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100010101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100010101101100) && ({row_reg, col_reg}<19'b0101100010101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100010101101111) && ({row_reg, col_reg}<19'b0101100010110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100010110010000) && ({row_reg, col_reg}<19'b0101100010110010010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0101100010110010010) && ({row_reg, col_reg}<19'b0101100010110010100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101100010110010100) && ({row_reg, col_reg}<19'b0101100010110011000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0101100010110011000) && ({row_reg, col_reg}<19'b0101100010110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100010110011101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101100010110011110)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101100010110011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101100010110100000) && ({row_reg, col_reg}<19'b0101100011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100011001010001) && ({row_reg, col_reg}<19'b0101100011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101100011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101100011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101100100000000000) && ({row_reg, col_reg}<19'b0101100100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100011110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101100100011110011) && ({row_reg, col_reg}<19'b0101100100011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100011111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101100100011111010) && ({row_reg, col_reg}<19'b0101100100011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100011111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101100100011111101) && ({row_reg, col_reg}<19'b0101100100100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100100100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100100100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101100100100000110) && ({row_reg, col_reg}<19'b0101100100100001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100100001000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101100100100001001) && ({row_reg, col_reg}<19'b0101100100100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100100100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100100100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101100100100010000) && ({row_reg, col_reg}<19'b0101100100100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101100100100010101) && ({row_reg, col_reg}<19'b0101100100100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0101100100100010111) && ({row_reg, col_reg}<19'b0101100100100011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100100100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100100100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100100100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100100100011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100100100011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101100100100100000) && ({row_reg, col_reg}<19'b0101100100100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100100100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100100100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100100100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100100100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100100110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100100100111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101100100100111001) && ({row_reg, col_reg}<19'b0101100100100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100100111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100100100111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101100100100111111) && ({row_reg, col_reg}<19'b0101100100101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100100101000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100100101000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100100101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100101001000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101100100101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100100101001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101100100101001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100100101001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100100101001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101100100101001110) && ({row_reg, col_reg}<19'b0101100100101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100101010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100100101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100101010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101100100101010100) && ({row_reg, col_reg}<19'b0101100100101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100100101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100101011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100100101011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100101011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101100100101011011) && ({row_reg, col_reg}<19'b0101100100101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100100101011110) && ({row_reg, col_reg}<19'b0101100100101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100101100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100101100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101100100101100011) && ({row_reg, col_reg}<19'b0101100100101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100101100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101100100101100111) && ({row_reg, col_reg}<19'b0101100100101101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100101101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101100100101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100100101101100) && ({row_reg, col_reg}<19'b0101100100101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100100101101111) && ({row_reg, col_reg}<19'b0101100100110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100110010000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0101100100110010001)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}>=19'b0101100100110010010) && ({row_reg, col_reg}<19'b0101100100110010100)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0101100100110010100) && ({row_reg, col_reg}<19'b0101100100110010110)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0101100100110010110) && ({row_reg, col_reg}<19'b0101100100110011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101100100110011000) && ({row_reg, col_reg}<19'b0101100100110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100100110011101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101100100110011110)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101100100110011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101100100110100000) && ({row_reg, col_reg}<19'b0101100101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100101001010001) && ({row_reg, col_reg}<19'b0101100101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101100101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101100101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101100110000000000) && ({row_reg, col_reg}<19'b0101100110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110011110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101100110011110011) && ({row_reg, col_reg}<19'b0101100110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110011111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100110011111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110011111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100110011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100110011111101) && ({row_reg, col_reg}<19'b0101100110011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100110100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100110100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100110100000110) && ({row_reg, col_reg}<19'b0101100110100001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110100001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101100110100001001) && ({row_reg, col_reg}<19'b0101100110100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100110100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100110100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101100110100010000) && ({row_reg, col_reg}<19'b0101100110100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101100110100010101) && ({row_reg, col_reg}<19'b0101100110100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110100010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101100110100011000) && ({row_reg, col_reg}<19'b0101100110100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100110100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110100011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101100110100011110) && ({row_reg, col_reg}<19'b0101100110100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100110100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100110100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101100110100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110100110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100110100111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101100110100111001) && ({row_reg, col_reg}<19'b0101100110100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110100111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100110100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110100111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100110100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100110101000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101100110101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101100110101000011) && ({row_reg, col_reg}<19'b0101100110101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110101000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101100110101000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100110101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110101001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100110101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100110101001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100110101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100110101001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100110101001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101100110101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100110101001111) && ({row_reg, col_reg}<19'b0101100110101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100110101010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100110101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110101010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100110101010100) && ({row_reg, col_reg}<19'b0101100110101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101100110101011000) && ({row_reg, col_reg}<19'b0101100110101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110101011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101100110101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101100110101011110) && ({row_reg, col_reg}<19'b0101100110101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110101100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101100110101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110101100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100110101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100110101100100) && ({row_reg, col_reg}<19'b0101100110101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101100110101100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100110101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110101101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101100110101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101100110101101100) && ({row_reg, col_reg}<19'b0101100110110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101100110110010000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101100110110010001) && ({row_reg, col_reg}<19'b0101100110110010011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0101100110110010011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0101100110110010100) && ({row_reg, col_reg}<19'b0101100110110010110)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0101100110110010110) && ({row_reg, col_reg}<19'b0101100110110011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101100110110011000) && ({row_reg, col_reg}<19'b0101100110110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100110110011101) && ({row_reg, col_reg}<19'b0101100110110100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101100110110100000) && ({row_reg, col_reg}<19'b0101100111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101100111001010001) && ({row_reg, col_reg}<19'b0101100111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101100111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101100111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101101000000000000) && ({row_reg, col_reg}<19'b0101101000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000011110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101101000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101101000011110011) && ({row_reg, col_reg}<19'b0101101000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000011111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101000011111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000011111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101000011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101000011111101) && ({row_reg, col_reg}<19'b0101101000011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101000100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101000100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101000100000110) && ({row_reg, col_reg}<19'b0101101000100001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101000100001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101101000100001001) && ({row_reg, col_reg}<19'b0101101000100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101000100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101000100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101000100010000) && ({row_reg, col_reg}<19'b0101101000100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101101000100010101) && ({row_reg, col_reg}<19'b0101101000100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000100010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101000100011000) && ({row_reg, col_reg}<19'b0101101000100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101000100011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101000100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000100011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101101000100011110) && ({row_reg, col_reg}<19'b0101101000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101000100101000) && ({row_reg, col_reg}<19'b0101101000100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101000100101101) && ({row_reg, col_reg}<19'b0101101000100110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101000100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101000100110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000100110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101000100111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101101000100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101000100111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101000100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000100111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101101000100111110) && ({row_reg, col_reg}<19'b0101101000101000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000101000110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101101000101000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101101000101001000) && ({row_reg, col_reg}<19'b0101101000101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000101001101) && ({row_reg, col_reg}<19'b0101101000101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101000101001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101101000101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101000101010001) && ({row_reg, col_reg}<19'b0101101000101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000101010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101101000101010100) && ({row_reg, col_reg}<19'b0101101000101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000101010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101101000101011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000101011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101000101011010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101101000101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101000101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101000101011110) && ({row_reg, col_reg}<19'b0101101000101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000101100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101101000101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000101100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101000101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101000101100100) && ({row_reg, col_reg}<19'b0101101000101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101000101100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101000101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000101101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101101000101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101000101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101000101101100) && ({row_reg, col_reg}<19'b0101101000110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101000110010000) && ({row_reg, col_reg}<19'b0101101000110010011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101101000110010011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0101101000110010100) && ({row_reg, col_reg}<19'b0101101000110011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101101000110011000) && ({row_reg, col_reg}<19'b0101101000110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101000110011101) && ({row_reg, col_reg}<19'b0101101000110100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101101000110100000) && ({row_reg, col_reg}<19'b0101101001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101001001010001) && ({row_reg, col_reg}<19'b0101101001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101101001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101101001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101101010000000000) && ({row_reg, col_reg}<19'b0101101010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010011110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101101010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101101010011110011) && ({row_reg, col_reg}<19'b0101101010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010011111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101101010011111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010011111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101010011111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101101010011111100) && ({row_reg, col_reg}<19'b0101101010011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101010011111110) && ({row_reg, col_reg}<19'b0101101010100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101010100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101010100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101010100000110) && ({row_reg, col_reg}<19'b0101101010100001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101010100001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101010100001001) && ({row_reg, col_reg}<19'b0101101010100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101010100001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101010100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101010100010000) && ({row_reg, col_reg}<19'b0101101010100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101010100010101) && ({row_reg, col_reg}<19'b0101101010100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010100010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101010100011000) && ({row_reg, col_reg}<19'b0101101010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101010100011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101010100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010100011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101010100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101010100100000) && ({row_reg, col_reg}<19'b0101101010100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101010100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101010100110110) && ({row_reg, col_reg}<19'b0101101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010100111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101101010100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101010100111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101101010100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010100111101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101101010100111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101010101000000) && ({row_reg, col_reg}<19'b0101101010101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101010101000010) && ({row_reg, col_reg}<19'b0101101010101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101010101000100) && ({row_reg, col_reg}<19'b0101101010101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010101000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101101010101001000) && ({row_reg, col_reg}<19'b0101101010101001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101010101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101010101001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101010101001101) && ({row_reg, col_reg}<19'b0101101010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010101001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101101010101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101010101010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010101010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101010101010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101010101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101010101010101) && ({row_reg, col_reg}<19'b0101101010101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101010101011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010101011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101101010101011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101010101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101010101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101010101011110) && ({row_reg, col_reg}<19'b0101101010101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010101100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101101010101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010101100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101010101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101010101100100) && ({row_reg, col_reg}<19'b0101101010101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101010101100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101010101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010101101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101101010101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101010101101100) && ({row_reg, col_reg}<19'b0101101010110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101010110001111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101101010110010000)) color_data = 12'b000000010011;
		if(({row_reg, col_reg}==19'b0101101010110010001)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}==19'b0101101010110010010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101101010110010011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101101010110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101010110010101) && ({row_reg, col_reg}<19'b0101101010110011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101101010110011000) && ({row_reg, col_reg}<19'b0101101010110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101010110011101) && ({row_reg, col_reg}<19'b0101101010110100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101101010110100000) && ({row_reg, col_reg}<19'b0101101011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101011001010001) && ({row_reg, col_reg}<19'b0101101011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101101011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101101011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101101100000000000) && ({row_reg, col_reg}<19'b0101101100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100011110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101101100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101101100011110011) && ({row_reg, col_reg}<19'b0101101100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100011111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101101100011111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100011111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101100011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101100011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100011111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101100011111110) && ({row_reg, col_reg}<19'b0101101100100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101100100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101100100000100) && ({row_reg, col_reg}<19'b0101101100100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100100000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101100100000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101100100001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101100100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101100100001010) && ({row_reg, col_reg}<19'b0101101100100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101100100001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101100100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101100100010000) && ({row_reg, col_reg}<19'b0101101100100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100100010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101100100010101) && ({row_reg, col_reg}<19'b0101101100100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100100010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101101100100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101100100011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101100100011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101100100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100100011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101100100011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101100100011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101100100100000) && ({row_reg, col_reg}<19'b0101101100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101100100110100) && ({row_reg, col_reg}<19'b0101101100100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100100110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101100100110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100100111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101101100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101100100111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101100100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101100100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101100100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101100101000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101100101000001) && ({row_reg, col_reg}<19'b0101101100101000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101100101000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101101100101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101100101000101) && ({row_reg, col_reg}<19'b0101101100101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100101000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101100101001000) && ({row_reg, col_reg}<19'b0101101100101001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101101100101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101100101001100) && ({row_reg, col_reg}<19'b0101101100101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101100101010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100101010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101100101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101100101010101) && ({row_reg, col_reg}<19'b0101101100101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100101010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101100101011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100101011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101100101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101100101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101100101011100) && ({row_reg, col_reg}<19'b0101101100101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101100101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101100101100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101100101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100101100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101101100101100011) && ({row_reg, col_reg}<19'b0101101100101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100101100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101101100101100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101100101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100101101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101101100101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101100101101100) && ({row_reg, col_reg}<19'b0101101100101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101100101101111) && ({row_reg, col_reg}<19'b0101101100110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101100110001010) && ({row_reg, col_reg}<19'b0101101100110010000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101101100110010000)) color_data = 12'b001101010111;
		if(({row_reg, col_reg}==19'b0101101100110010001)) color_data = 12'b001001000110;
		if(({row_reg, col_reg}==19'b0101101100110010010)) color_data = 12'b000000100100;
		if(({row_reg, col_reg}==19'b0101101100110010011)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}>=19'b0101101100110010100) && ({row_reg, col_reg}<19'b0101101100110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101100110010110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0101101100110010111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0101101100110011000) && ({row_reg, col_reg}<19'b0101101100110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101100110011101) && ({row_reg, col_reg}<19'b0101101100110100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101101100110100000) && ({row_reg, col_reg}<19'b0101101101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101101001010001) && ({row_reg, col_reg}<19'b0101101101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101101101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101101101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101101110000000000) && ({row_reg, col_reg}<19'b0101101110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110011110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101101110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101101110011110011) && ({row_reg, col_reg}<19'b0101101110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101110011111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110011111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101101110011111011) && ({row_reg, col_reg}<19'b0101101110011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110011111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101110100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110100000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101110100000100) && ({row_reg, col_reg}<19'b0101101110100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101110100000110) && ({row_reg, col_reg}<19'b0101101110100001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101110100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101110100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101110100001010) && ({row_reg, col_reg}<19'b0101101110100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101110100001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101110100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101110100010000) && ({row_reg, col_reg}<19'b0101101110100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110100010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101110100010101) && ({row_reg, col_reg}<19'b0101101110100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110100010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101101110100011000) && ({row_reg, col_reg}<19'b0101101110100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110100011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101101110100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110100011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101101110100011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101110100011111) && ({row_reg, col_reg}<19'b0101101110100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101110100110100) && ({row_reg, col_reg}<19'b0101101110100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110100110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101110100110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101101110100111001) && ({row_reg, col_reg}<19'b0101101110100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110100111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101110100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110100111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101110100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101110101000001) && ({row_reg, col_reg}<19'b0101101110101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101110101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101110101000101) && ({row_reg, col_reg}<19'b0101101110101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101110101001000) && ({row_reg, col_reg}<19'b0101101110101001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101110101001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101101110101001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101110101001111) && ({row_reg, col_reg}<19'b0101101110101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110101010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101110101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101110101010101) && ({row_reg, col_reg}<19'b0101101110101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101110101011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101110101011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101110101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101110101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101110101011100) && ({row_reg, col_reg}<19'b0101101110101011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101101110101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101101110101100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101110101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110101100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101101110101100011) && ({row_reg, col_reg}<19'b0101101110101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101101110101100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101110101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110101101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101101110101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101101110101101100) && ({row_reg, col_reg}<19'b0101101110101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101101110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101101110101101111) && ({row_reg, col_reg}<19'b0101101110110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101110110001000) && ({row_reg, col_reg}<19'b0101101110110001101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101101110110001101) && ({row_reg, col_reg}<19'b0101101110110010000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101101110110010000)) color_data = 12'b011110001100;
		if(({row_reg, col_reg}==19'b0101101110110010001)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==19'b0101101110110010010)) color_data = 12'b001001000111;
		if(({row_reg, col_reg}==19'b0101101110110010011)) color_data = 12'b000000010011;
		if(({row_reg, col_reg}==19'b0101101110110010100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101101110110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101110110010110) && ({row_reg, col_reg}<19'b0101101110110011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101101110110011000) && ({row_reg, col_reg}<19'b0101101110110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101110110011110) && ({row_reg, col_reg}<19'b0101101110110100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101101110110100000) && ({row_reg, col_reg}<19'b0101101111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101101111001010001) && ({row_reg, col_reg}<19'b0101101111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101101111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101101111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101110000000000000) && ({row_reg, col_reg}<19'b0101110000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101110000011110011) && ({row_reg, col_reg}<19'b0101110000011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000011111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110000011111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000011111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101110000011111011) && ({row_reg, col_reg}<19'b0101110000011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110000011111110) && ({row_reg, col_reg}<19'b0101110000100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110000100000100) && ({row_reg, col_reg}<19'b0101110000100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110000100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110000100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110000100001010) && ({row_reg, col_reg}<19'b0101110000100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110000100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110000100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110000100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101110000100010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000100010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110000100010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101110000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110000100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110000100011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110000100011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101110000100100000) && ({row_reg, col_reg}<19'b0101110000100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110000100100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110000100100110) && ({row_reg, col_reg}<19'b0101110000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110000100101001) && ({row_reg, col_reg}<19'b0101110000100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110000100101011) && ({row_reg, col_reg}<19'b0101110000100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110000100101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101110000100110000) && ({row_reg, col_reg}<19'b0101110000100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110000100110100) && ({row_reg, col_reg}<19'b0101110000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110000100110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000100111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110000100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110000100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000100111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110000100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000100111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110000100111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110000101000000) && ({row_reg, col_reg}<19'b0101110000101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000101010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101110000101010001) && ({row_reg, col_reg}<19'b0101110000101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000101010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101110000101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110000101010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110000101011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110000101011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110000101011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000101011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110000101011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101110000101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110000101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000101100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110000101100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110000101100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101110000101100011) && ({row_reg, col_reg}<19'b0101110000101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110000101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110000101100111) && ({row_reg, col_reg}<19'b0101110000101101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000101101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110000101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101110000101101100) && ({row_reg, col_reg}<19'b0101110000110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110000110000111) && ({row_reg, col_reg}<19'b0101110000110001001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110000110001001)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0101110000110001010) && ({row_reg, col_reg}<19'b0101110000110001100)) color_data = 12'b000100010011;
		if(({row_reg, col_reg}==19'b0101110000110001100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}>=19'b0101110000110001101) && ({row_reg, col_reg}<19'b0101110000110001111)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101110000110001111)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101110000110010000)) color_data = 12'b011001111011;
		if(({row_reg, col_reg}==19'b0101110000110010001)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==19'b0101110000110010010)) color_data = 12'b001001000111;
		if(({row_reg, col_reg}==19'b0101110000110010011)) color_data = 12'b000000100101;
		if(({row_reg, col_reg}==19'b0101110000110010100)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}==19'b0101110000110010101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110000110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110000110010111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101110000110011000) && ({row_reg, col_reg}<19'b0101110000110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110000110011110) && ({row_reg, col_reg}<19'b0101110000110100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101110000110100000) && ({row_reg, col_reg}<19'b0101110001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110001001010001) && ({row_reg, col_reg}<19'b0101110001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101110001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101110010000000000) && ({row_reg, col_reg}<19'b0101110010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101110010011110011) && ({row_reg, col_reg}<19'b0101110010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010011111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110010011111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010011111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101110010011111011) && ({row_reg, col_reg}<19'b0101110010011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110010011111110) && ({row_reg, col_reg}<19'b0101110010100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110010100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110010100000100) && ({row_reg, col_reg}<19'b0101110010100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110010100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101110010100001001) && ({row_reg, col_reg}<19'b0101110010100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110010100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110010100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110010100010001) && ({row_reg, col_reg}<19'b0101110010100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110010100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101110010100010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110010100010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110010100010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110010100011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110010100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010100011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110010100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101110010100100001) && ({row_reg, col_reg}<19'b0101110010100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110010100100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110010100101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101110010100101001) && ({row_reg, col_reg}<19'b0101110010100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110010100110100) && ({row_reg, col_reg}<19'b0101110010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110010100110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010100111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110010100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110010100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010100111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110010100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010100111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110010100111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101110010100111111) && ({row_reg, col_reg}<19'b0101110010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110010101010001) && ({row_reg, col_reg}<19'b0101110010101010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110010101010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101110010101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110010101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110010101010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110010101011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110010101011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101110010101011010) && ({row_reg, col_reg}<19'b0101110010101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010101011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110010101011101) && ({row_reg, col_reg}<19'b0101110010101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010101011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110010101100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110010101100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110010101100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101110010101100011) && ({row_reg, col_reg}<19'b0101110010101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110010101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110010101100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010101101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110010101101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110010101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101110010101101100) && ({row_reg, col_reg}<19'b0101110010101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110010101101111) && ({row_reg, col_reg}<19'b0101110010110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010110000111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101110010110001000) && ({row_reg, col_reg}<19'b0101110010110001010)) color_data = 12'b000100010011;
		if(({row_reg, col_reg}==19'b0101110010110001010)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}>=19'b0101110010110001011) && ({row_reg, col_reg}<19'b0101110010110001110)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101110010110001110)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==19'b0101110010110001111)) color_data = 12'b001000100111;
		if(({row_reg, col_reg}==19'b0101110010110010000)) color_data = 12'b011001111100;
		if(({row_reg, col_reg}==19'b0101110010110010001)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==19'b0101110010110010010)) color_data = 12'b001001001000;
		if(({row_reg, col_reg}==19'b0101110010110010011)) color_data = 12'b000000100101;
		if(({row_reg, col_reg}==19'b0101110010110010100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101110010110010101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110010110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110010110010111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101110010110011000) && ({row_reg, col_reg}<19'b0101110010110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110010110011110) && ({row_reg, col_reg}<19'b0101110010110100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101110010110100000) && ({row_reg, col_reg}<19'b0101110011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110011001010001) && ({row_reg, col_reg}<19'b0101110011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101110011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101110100000000000) && ({row_reg, col_reg}<19'b0101110100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101110100011110011) && ({row_reg, col_reg}<19'b0101110100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100011111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110100011111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100011111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101110100011111011) && ({row_reg, col_reg}<19'b0101110100011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110100011111110) && ({row_reg, col_reg}<19'b0101110100100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110100100000100) && ({row_reg, col_reg}<19'b0101110100100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110100100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101110100100001001) && ({row_reg, col_reg}<19'b0101110100100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110100100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110100100010001) && ({row_reg, col_reg}<19'b0101110100100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100100010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110100100010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100100010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110100100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110100100011010) && ({row_reg, col_reg}<19'b0101110100100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100100011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101110100100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110100100011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110100100100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110100100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110100100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110100100100011) && ({row_reg, col_reg}<19'b0101110100100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110100100100101) && ({row_reg, col_reg}<19'b0101110100100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110100100101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110100100101010) && ({row_reg, col_reg}<19'b0101110100100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110100100101111) && ({row_reg, col_reg}<19'b0101110100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110100100110100) && ({row_reg, col_reg}<19'b0101110100100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100100110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110100100111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100100111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110100100111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101110100100111111) && ({row_reg, col_reg}<19'b0101110100101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100101010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110100101010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110100101010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110100101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100101010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110100101011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110100101011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110100101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110100101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110100101011100) && ({row_reg, col_reg}<19'b0101110100101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110100101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100101100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110100101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100101100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101110100101100011) && ({row_reg, col_reg}<19'b0101110100101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110100101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100101100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100101100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110100101101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110100101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110100101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101110100101101100) && ({row_reg, col_reg}<19'b0101110100101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110100101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110100101101111) && ({row_reg, col_reg}<19'b0101110100110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110100110000110) && ({row_reg, col_reg}<19'b0101110100110001000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110100110001000)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0101110100110001001)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}>=19'b0101110100110001010) && ({row_reg, col_reg}<19'b0101110100110001101)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101110100110001101)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0101110100110001110)) color_data = 12'b001100100111;
		if(({row_reg, col_reg}==19'b0101110100110001111)) color_data = 12'b010101011010;
		if(({row_reg, col_reg}==19'b0101110100110010000)) color_data = 12'b011001111101;
		if(({row_reg, col_reg}==19'b0101110100110010001)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==19'b0101110100110010010)) color_data = 12'b000100111000;
		if(({row_reg, col_reg}==19'b0101110100110010011)) color_data = 12'b000000010101;
		if(({row_reg, col_reg}==19'b0101110100110010100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0101110100110010101) && ({row_reg, col_reg}<19'b0101110100110010111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110100110010111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0101110100110011000) && ({row_reg, col_reg}<19'b0101110101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110101001010001) && ({row_reg, col_reg}<19'b0101110101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101110101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101110110000000000) && ({row_reg, col_reg}<19'b0101110110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101110110011110011) && ({row_reg, col_reg}<19'b0101110110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110011111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110110011111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110011111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101110110011111011) && ({row_reg, col_reg}<19'b0101110110100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110110100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110110100000100) && ({row_reg, col_reg}<19'b0101110110100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110110100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101110110100001001) && ({row_reg, col_reg}<19'b0101110110100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110110100001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110110100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110110100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110110100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110110100010001) && ({row_reg, col_reg}<19'b0101110110100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101110110100010011) && ({row_reg, col_reg}<19'b0101110110100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110100010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110110100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110100011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101110110100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110110100011011) && ({row_reg, col_reg}<19'b0101110110100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110110100011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110110100011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110100011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110110100100001) && ({row_reg, col_reg}<19'b0101110110100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110110100100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101110110100100101) && ({row_reg, col_reg}<19'b0101110110100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110110100101011) && ({row_reg, col_reg}<19'b0101110110100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110110100101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110110100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110110100110000) && ({row_reg, col_reg}<19'b0101110110100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110110100110100) && ({row_reg, col_reg}<19'b0101110110100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101110110100110111) && ({row_reg, col_reg}<19'b0101110110100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110100111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101110110100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110100111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101110110100111100) && ({row_reg, col_reg}<19'b0101110110100111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110110100111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101110110100111111) && ({row_reg, col_reg}<19'b0101110110101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110101010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110110101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110101010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110110101010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110110101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110110101010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110110101011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110101011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110110101011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110110101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110101011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101110110101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110110101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101110110101100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101110110101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101110110101100011) && ({row_reg, col_reg}<19'b0101110110101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110110101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110101100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101110110101100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110101101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110110101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101110110101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110110101101100) && ({row_reg, col_reg}<19'b0101110110101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101110110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101110110101101111) && ({row_reg, col_reg}<19'b0101110110110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110110110000110) && ({row_reg, col_reg}<19'b0101110110110001000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110110110001000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0101110110110001001) && ({row_reg, col_reg}<19'b0101110110110001100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101110110110001100)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0101110110110001101)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==19'b0101110110110001110)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==19'b0101110110110001111)) color_data = 12'b011001011011;
		if(({row_reg, col_reg}==19'b0101110110110010000)) color_data = 12'b011001111101;
		if(({row_reg, col_reg}==19'b0101110110110010001)) color_data = 12'b010001011100;
		if(({row_reg, col_reg}==19'b0101110110110010010)) color_data = 12'b001000111001;
		if(({row_reg, col_reg}==19'b0101110110110010011)) color_data = 12'b000000010110;
		if(({row_reg, col_reg}==19'b0101110110110010100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101110110110010101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101110110110010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110110110010111)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0101110110110011000) && ({row_reg, col_reg}<19'b0101110111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101110111001010001) && ({row_reg, col_reg}<19'b0101110111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101110111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101110111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101111000000000000) && ({row_reg, col_reg}<19'b0101111000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101111000011110011) && ({row_reg, col_reg}<19'b0101111000011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000011111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111000011111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000011111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111000011111011) && ({row_reg, col_reg}<19'b0101111000011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111000100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111000100000100) && ({row_reg, col_reg}<19'b0101111000100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111000100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000100001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101111000100001001) && ({row_reg, col_reg}<19'b0101111000100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111000100001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101111000100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111000100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111000100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111000100010001) && ({row_reg, col_reg}<19'b0101111000100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111000100010011) && ({row_reg, col_reg}<19'b0101111000100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101111000100010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111000100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000100011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101111000100011001) && ({row_reg, col_reg}<19'b0101111000100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111000100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101111000100011110) && ({row_reg, col_reg}<19'b0101111000100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000100100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101111000100100001) && ({row_reg, col_reg}<19'b0101111000100100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111000100100101) && ({row_reg, col_reg}<19'b0101111000100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101111000100101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000100101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101111000100101100) && ({row_reg, col_reg}<19'b0101111000100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111000100110100) && ({row_reg, col_reg}<19'b0101111000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101111000100110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000100111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101111000100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111000100111100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111000100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111000100111111) && ({row_reg, col_reg}<19'b0101111000101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111000101010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101111000101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111000101010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101111000101011000) && ({row_reg, col_reg}<19'b0101111000101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000101011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101111000101011011) && ({row_reg, col_reg}<19'b0101111000101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111000101011101) && ({row_reg, col_reg}<19'b0101111000101011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111000101011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101111000101100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000101100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111000101100010) && ({row_reg, col_reg}<19'b0101111000101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111000101100110) && ({row_reg, col_reg}<19'b0101111000101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101111000101101001) && ({row_reg, col_reg}<19'b0101111000101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111000101101100) && ({row_reg, col_reg}<19'b0101111000101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111000101101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111000101101111) && ({row_reg, col_reg}<19'b0101111000110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111000110000110) && ({row_reg, col_reg}<19'b0101111000110001000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101111000110001000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101111000110001001)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101111000110001010)) color_data = 12'b000100010101;
		if(({row_reg, col_reg}==19'b0101111000110001011)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==19'b0101111000110001100)) color_data = 12'b001000010111;
		if(({row_reg, col_reg}==19'b0101111000110001101)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==19'b0101111000110001110)) color_data = 12'b010101001010;
		if(({row_reg, col_reg}==19'b0101111000110001111)) color_data = 12'b011001101100;
		if(({row_reg, col_reg}==19'b0101111000110010000)) color_data = 12'b011001101110;
		if(({row_reg, col_reg}==19'b0101111000110010001)) color_data = 12'b010001101101;
		if(({row_reg, col_reg}==19'b0101111000110010010)) color_data = 12'b001001001010;
		if(({row_reg, col_reg}==19'b0101111000110010011)) color_data = 12'b000000100111;
		if(({row_reg, col_reg}==19'b0101111000110010100)) color_data = 12'b000000010101;
		if(({row_reg, col_reg}==19'b0101111000110010101)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}>=19'b0101111000110010110) && ({row_reg, col_reg}<19'b0101111000110011000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0101111000110011000) && ({row_reg, col_reg}<19'b0101111001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111001001010001) && ({row_reg, col_reg}<19'b0101111001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101111001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101111001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101111010000000000) && ({row_reg, col_reg}<19'b0101111010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101111010011110011) && ({row_reg, col_reg}<19'b0101111010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010011111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111010011111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111010011111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111010011111011) && ({row_reg, col_reg}<19'b0101111010011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111010100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111010100000100) && ({row_reg, col_reg}<19'b0101111010100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111010100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010100001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101111010100001001) && ({row_reg, col_reg}<19'b0101111010100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111010100001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101111010100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111010100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111010100010001) && ({row_reg, col_reg}<19'b0101111010100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111010100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111010100010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111010100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111010100011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111010100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111010100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111010100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111010100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010100100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111010100100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101111010100100010) && ({row_reg, col_reg}<19'b0101111010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111010100100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101111010100100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111010100101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111010100101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111010100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010100101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111010100101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101111010100101101) && ({row_reg, col_reg}<19'b0101111010100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111010100110100) && ({row_reg, col_reg}<19'b0101111010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101111010100110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010100111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111010100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010100111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111010100111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111010100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010100111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111010100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111010101000000) && ({row_reg, col_reg}<19'b0101111010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111010101010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101111010101010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111010101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010101010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101111010101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111010101010110) && ({row_reg, col_reg}<19'b0101111010101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111010101011000) && ({row_reg, col_reg}<19'b0101111010101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010101011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101111010101011011) && ({row_reg, col_reg}<19'b0101111010101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010101011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101111010101011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111010101100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111010101100010) && ({row_reg, col_reg}<19'b0101111010101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010101100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101111010101100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010101100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111010101101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101111010101101001) && ({row_reg, col_reg}<19'b0101111010101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111010101101100) && ({row_reg, col_reg}<19'b0101111010101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010101101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111010101101111) && ({row_reg, col_reg}<19'b0101111010110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111010110000110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101111010110000111)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101111010110001000)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101111010110001001)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==19'b0101111010110001010)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==19'b0101111010110001011)) color_data = 12'b010101011010;
		if(({row_reg, col_reg}==19'b0101111010110001100)) color_data = 12'b011001011011;
		if(({row_reg, col_reg}==19'b0101111010110001101)) color_data = 12'b011001011100;
		if(({row_reg, col_reg}==19'b0101111010110001110)) color_data = 12'b011101101100;
		if(({row_reg, col_reg}==19'b0101111010110001111)) color_data = 12'b011101111110;
		if(({row_reg, col_reg}==19'b0101111010110010000)) color_data = 12'b010101101110;
		if(({row_reg, col_reg}==19'b0101111010110010001)) color_data = 12'b010001101101;
		if(({row_reg, col_reg}==19'b0101111010110010010)) color_data = 12'b001101011100;
		if(({row_reg, col_reg}==19'b0101111010110010011)) color_data = 12'b001001001001;
		if(({row_reg, col_reg}==19'b0101111010110010100)) color_data = 12'b000100110111;
		if(({row_reg, col_reg}==19'b0101111010110010101)) color_data = 12'b000000010100;
		if(({row_reg, col_reg}==19'b0101111010110010110)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0101111010110010111) && ({row_reg, col_reg}<19'b0101111011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111011001010001) && ({row_reg, col_reg}<19'b0101111011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101111011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101111011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101111100000000000) && ({row_reg, col_reg}<19'b0101111100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101111100011110011) && ({row_reg, col_reg}<19'b0101111100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111100011111000) && ({row_reg, col_reg}<19'b0101111100011111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111100011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101111100011111011) && ({row_reg, col_reg}<19'b0101111100011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111100100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111100100000100) && ({row_reg, col_reg}<19'b0101111100100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111100100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100100001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101111100100001001) && ({row_reg, col_reg}<19'b0101111100100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111100100001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101111100100001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111100100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111100100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111100100010001) && ({row_reg, col_reg}<19'b0101111100100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111100100010100) && ({row_reg, col_reg}<19'b0101111100100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101111100100010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111100100011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111100100011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111100100011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111100100011011) && ({row_reg, col_reg}<19'b0101111100100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101111100100011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111100100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100100100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101111100100100010) && ({row_reg, col_reg}<19'b0101111100100100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101111100100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111100100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111100100100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101111100100100111) && ({row_reg, col_reg}<19'b0101111100100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0101111100100101001) && ({row_reg, col_reg}<19'b0101111100100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111100100101011) && ({row_reg, col_reg}<19'b0101111100100101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100100101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0101111100100101110) && ({row_reg, col_reg}<19'b0101111100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111100100110100) && ({row_reg, col_reg}<19'b0101111100100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101111100100110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100100111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111100100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111100100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111100100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111100100111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111100101000000) && ({row_reg, col_reg}<19'b0101111100101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111100101010000) && ({row_reg, col_reg}<19'b0101111100101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111100101010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111100101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100101010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101111100101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111100101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111100101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111100101011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100101011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111100101011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101111100101011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0101111100101011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0101111100101011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111100101011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100101100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111100101100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111100101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111100101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111100101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100101100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111100101100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111100101100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111100101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111100101101001) && ({row_reg, col_reg}<19'b0101111100101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111100101101100) && ({row_reg, col_reg}<19'b0101111100101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100101101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111100101101111) && ({row_reg, col_reg}<19'b0101111100110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111100110000110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101111100110000111)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101111100110001000)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0101111100110001001)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==19'b0101111100110001010)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==19'b0101111100110001011)) color_data = 12'b011001011010;
		if(({row_reg, col_reg}==19'b0101111100110001100)) color_data = 12'b011001011011;
		if(({row_reg, col_reg}==19'b0101111100110001101)) color_data = 12'b011001011100;
		if(({row_reg, col_reg}==19'b0101111100110001110)) color_data = 12'b011101101101;
		if(({row_reg, col_reg}==19'b0101111100110001111)) color_data = 12'b011101111110;
		if(({row_reg, col_reg}==19'b0101111100110010000)) color_data = 12'b010101011110;
		if(({row_reg, col_reg}==19'b0101111100110010001)) color_data = 12'b010001101110;
		if(({row_reg, col_reg}==19'b0101111100110010010)) color_data = 12'b010101101101;
		if(({row_reg, col_reg}==19'b0101111100110010011)) color_data = 12'b010001101100;
		if(({row_reg, col_reg}==19'b0101111100110010100)) color_data = 12'b001101011001;
		if(({row_reg, col_reg}==19'b0101111100110010101)) color_data = 12'b000100110110;
		if(({row_reg, col_reg}==19'b0101111100110010110)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}>=19'b0101111100110010111) && ({row_reg, col_reg}<19'b0101111101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111101001010001) && ({row_reg, col_reg}<19'b0101111101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101111101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101111101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0101111110000000000) && ({row_reg, col_reg}<19'b0101111110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111110011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101111110011110011) && ({row_reg, col_reg}<19'b0101111110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111110011111000) && ({row_reg, col_reg}<19'b0101111110011111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111110011111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101111110011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110011111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111110011111101) && ({row_reg, col_reg}<19'b0101111110011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111110100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111110100000100) && ({row_reg, col_reg}<19'b0101111110100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111110100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110100001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101111110100001001) && ({row_reg, col_reg}<19'b0101111110100001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111110100001100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101111110100001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111110100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0101111110100001111) && ({row_reg, col_reg}<19'b0101111110100010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111110100010001) && ({row_reg, col_reg}<19'b0101111110100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111110100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111110100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111110100010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111110100011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111110100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110100011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101111110100011011) && ({row_reg, col_reg}<19'b0101111110100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0101111110100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101111110100100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111110100100011) && ({row_reg, col_reg}<19'b0101111110100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111110100101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111110100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101111110100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111110100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110100101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0101111110100101110) && ({row_reg, col_reg}<19'b0101111110100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0101111110100110100) && ({row_reg, col_reg}<19'b0101111110100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0101111110100110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110100111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111110100111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111110100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111110100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110100111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111110100111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101111110101000000) && ({row_reg, col_reg}<19'b0101111110101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111110101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111110101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111110101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111110101010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101111110101010111) && ({row_reg, col_reg}<19'b0101111110101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110101011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111110101011010) && ({row_reg, col_reg}<19'b0101111110101011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110101011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101111110101011101) && ({row_reg, col_reg}<19'b0101111110101011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111110101011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110101100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111110101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110101100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0101111110101100011) && ({row_reg, col_reg}<19'b0101111110101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0101111110101100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101111110101100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111110101100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111110101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0101111110101101001) && ({row_reg, col_reg}<19'b0101111110101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110101101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111110101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0101111110101101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0101111110101101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0101111110101101111) && ({row_reg, col_reg}<19'b0101111110110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111110110000110) && ({row_reg, col_reg}<19'b0101111110110001000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101111110110001000)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0101111110110001001)) color_data = 12'b000100010100;
		if(({row_reg, col_reg}==19'b0101111110110001010)) color_data = 12'b001100100110;
		if(({row_reg, col_reg}==19'b0101111110110001011)) color_data = 12'b001100110111;
		if(({row_reg, col_reg}==19'b0101111110110001100)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==19'b0101111110110001101)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}==19'b0101111110110001110)) color_data = 12'b010101011010;
		if(({row_reg, col_reg}==19'b0101111110110001111)) color_data = 12'b011001101100;
		if(({row_reg, col_reg}==19'b0101111110110010000)) color_data = 12'b010101011100;
		if(({row_reg, col_reg}==19'b0101111110110010001)) color_data = 12'b010101101101;
		if(({row_reg, col_reg}==19'b0101111110110010010)) color_data = 12'b011001111101;
		if(({row_reg, col_reg}==19'b0101111110110010011)) color_data = 12'b011001111100;
		if(({row_reg, col_reg}==19'b0101111110110010100)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==19'b0101111110110010101)) color_data = 12'b001000110110;
		if(({row_reg, col_reg}==19'b0101111110110010110)) color_data = 12'b000000010010;
		if(({row_reg, col_reg}>=19'b0101111110110010111) && ({row_reg, col_reg}<19'b0101111111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0101111111001010001) && ({row_reg, col_reg}<19'b0101111111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0101111111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0101111111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110000000000000000) && ({row_reg, col_reg}<19'b0110000000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000011110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000011110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000000011110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110000000011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000000011110101) && ({row_reg, col_reg}<19'b0110000000011110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000000011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000011111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000000011111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000000011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000000011111100) && ({row_reg, col_reg}<19'b0110000000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000000011111111) && ({row_reg, col_reg}<19'b0110000000100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000000100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000000100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000100001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000000100001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110000000100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000100001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000000100001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000000100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000100001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000000100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110000000100010000) && ({row_reg, col_reg}<19'b0110000000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000000100011000) && ({row_reg, col_reg}<19'b0110000000100011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000000100011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000000100011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000000100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000000100011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000000100011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000000100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000000100100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000000100100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000000100100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000000100100100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000000100100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000000100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000000100100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110000000100101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000000100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000000100101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000100101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0110000000100101110) && ({row_reg, col_reg}<19'b0110000000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000000100110110) && ({row_reg, col_reg}<19'b0110000000100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000100111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000000100111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110000000100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000000100111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000000100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000100111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110000000101000000) && ({row_reg, col_reg}<19'b0110000000101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000101010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000000101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000101010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000000101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000000101010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110000000101010110) && ({row_reg, col_reg}<19'b0110000000101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000101011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000000101011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0110000000101011011) && ({row_reg, col_reg}<19'b0110000000101011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000101011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000000101011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000000101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000101100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110000000101100010) && ({row_reg, col_reg}<19'b0110000000101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000101100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110000000101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000101100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110000000101100111) && ({row_reg, col_reg}<19'b0110000000110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000000110001000)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b0110000000110001001) && ({row_reg, col_reg}<19'b0110000000110001110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110000000110001110)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==19'b0110000000110001111)) color_data = 12'b011001101001;
		if(({row_reg, col_reg}>=19'b0110000000110010000) && ({row_reg, col_reg}<19'b0110000000110010010)) color_data = 12'b011001101011;
		if(({row_reg, col_reg}==19'b0110000000110010010)) color_data = 12'b011001011010;
		if(({row_reg, col_reg}==19'b0110000000110010011)) color_data = 12'b010001001000;
		if(({row_reg, col_reg}==19'b0110000000110010100)) color_data = 12'b000100010101;
		if(({row_reg, col_reg}==19'b0110000000110010101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0110000000110010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110000000110010111) && ({row_reg, col_reg}<19'b0110000001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000001001010001) && ({row_reg, col_reg}<19'b0110000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110000001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110000001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110000010000000000) && ({row_reg, col_reg}<19'b0110000010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010011110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000010011110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000010011110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000010011110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0110000010011110100) && ({row_reg, col_reg}<19'b0110000010011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000010011110110) && ({row_reg, col_reg}<19'b0110000010011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000010011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010011111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000010011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0110000010011111011) && ({row_reg, col_reg}<19'b0110000010011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000010011111101) && ({row_reg, col_reg}<19'b0110000010011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000010011111111) && ({row_reg, col_reg}<19'b0110000010100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000010100000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000010100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010100001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000010100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110000010100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010100001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000010100001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000010100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010100001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000010100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000010100010000) && ({row_reg, col_reg}<19'b0110000010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010100011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110000010100011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000010100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010100011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0110000010100011100) && ({row_reg, col_reg}<19'b0110000010100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010100011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000010100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000010100100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000010100100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000010100100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000010100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000010100100110) && ({row_reg, col_reg}<19'b0110000010100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010100101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110000010100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010100101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000010100101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000010100110000) && ({row_reg, col_reg}<19'b0110000010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000010100110110) && ({row_reg, col_reg}<19'b0110000010100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010100111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000010100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000010100111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010100111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000010100111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000010100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010100111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110000010101000000) && ({row_reg, col_reg}<19'b0110000010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000010101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010101010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000010101010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000010101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010101010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000010101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110000010101010111) && ({row_reg, col_reg}<19'b0110000010101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000010101011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000010101011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110000010101011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110000010101011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110000010101011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110000010101011111) && ({row_reg, col_reg}<19'b0110000010101100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110000010101100001) && ({row_reg, col_reg}<19'b0110000010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010101100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110000010101100100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000010101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010101100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000010101100111) && ({row_reg, col_reg}<19'b0110000010110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010110001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110000010110001001) && ({row_reg, col_reg}<19'b0110000010110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000010110001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000010110001111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==19'b0110000010110010000)) color_data = 12'b011001011000;
		if(({row_reg, col_reg}==19'b0110000010110010001)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==19'b0110000010110010010)) color_data = 12'b001100110111;
		if(({row_reg, col_reg}==19'b0110000010110010011)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==19'b0110000010110010100)) color_data = 12'b000100010011;
		if(({row_reg, col_reg}==19'b0110000010110010101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0110000010110010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110000010110010111) && ({row_reg, col_reg}<19'b0110000011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000011001010001) && ({row_reg, col_reg}<19'b0110000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110000011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110000011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110000100000000000) && ({row_reg, col_reg}<19'b0110000100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100011110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110000100011110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000100011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100011110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0110000100011110100) && ({row_reg, col_reg}<19'b0110000100011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100011110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000100011110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110000100011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100011111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000100011111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0110000100011111011) && ({row_reg, col_reg}<19'b0110000100011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000100011111101) && ({row_reg, col_reg}<19'b0110000100011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000100011111111) && ({row_reg, col_reg}<19'b0110000100100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000100100000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000100100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000100100001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000100100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100100001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110000100100001100) && ({row_reg, col_reg}<19'b0110000100100001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000100100001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0110000100100001111) && ({row_reg, col_reg}<19'b0110000100100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100100011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0110000100100011010) && ({row_reg, col_reg}<19'b0110000100100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100100011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0110000100100011101) && ({row_reg, col_reg}<19'b0110000100100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100100101001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110000100100101010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000100100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100100101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000100100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000100100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000100100110000) && ({row_reg, col_reg}<19'b0110000100100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000100100110110) && ({row_reg, col_reg}<19'b0110000100100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000100100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000100100111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000100100111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0110000100100111011) && ({row_reg, col_reg}<19'b0110000100100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100100111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000100100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100100111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0110000100101000000) && ({row_reg, col_reg}<19'b0110000100101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000100101010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000100101010100) && ({row_reg, col_reg}<19'b0110000100101010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100101010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000100101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110000100101011001) && ({row_reg, col_reg}<19'b0110000100101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100101100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000100101100001) && ({row_reg, col_reg}<19'b0110000100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100101100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000100101100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100101100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000100101100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110000100101100111) && ({row_reg, col_reg}<19'b0110000100110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000100110001001) && ({row_reg, col_reg}<19'b0110000100110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000100110001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000100110001111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==19'b0110000100110010000)) color_data = 12'b010101011000;
		if(({row_reg, col_reg}==19'b0110000100110010001)) color_data = 12'b001100100110;
		if(({row_reg, col_reg}==19'b0110000100110010010)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==19'b0110000100110010011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0110000100110010100)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==19'b0110000100110010101)) color_data = 12'b000100010011;
		if(({row_reg, col_reg}==19'b0110000100110010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110000100110010111) && ({row_reg, col_reg}<19'b0110000101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000101001010001) && ({row_reg, col_reg}<19'b0110000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110000101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110000101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110000110000000000) && ({row_reg, col_reg}<19'b0110000110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110011110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000110011110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000110011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110011110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0110000110011110100) && ({row_reg, col_reg}<19'b0110000110011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110011110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000110011110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110000110011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110011111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000110011111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110000110011111011) && ({row_reg, col_reg}<19'b0110000110011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000110011111101) && ({row_reg, col_reg}<19'b0110000110011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000110011111111) && ({row_reg, col_reg}<19'b0110000110100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000110100000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110000110100000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000110100001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000110100001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000110100001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110000110100001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000110100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110100001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000110100001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110000110100001111) && ({row_reg, col_reg}<19'b0110000110100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110100011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000110100011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000110100011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000110100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110100011101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000110100011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110000110100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110100100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000110100100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000110100100010) && ({row_reg, col_reg}<19'b0110000110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000110100100110) && ({row_reg, col_reg}<19'b0110000110100101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000110100101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000110100101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110000110100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110100101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000110100101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110000110100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000110100101110) && ({row_reg, col_reg}<19'b0110000110100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110000110100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0110000110100111001) && ({row_reg, col_reg}<19'b0110000110100111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000110100111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000110100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110100111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000110100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0110000110101000000) && ({row_reg, col_reg}<19'b0110000110101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110101010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000110101010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000110101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110101010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110000110101010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110000110101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000110101011001) && ({row_reg, col_reg}<19'b0110000110101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110101011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110000110101011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000110101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000110101011111) && ({row_reg, col_reg}<19'b0110000110101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110101100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110000110101100011) && ({row_reg, col_reg}<19'b0110000110101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110101100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110000110101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110000110101101000) && ({row_reg, col_reg}<19'b0110000110110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110000110110001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110000110110001111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==19'b0110000110110010000)) color_data = 12'b011001101001;
		if(({row_reg, col_reg}==19'b0110000110110010001)) color_data = 12'b001100100110;
		if(({row_reg, col_reg}>=19'b0110000110110010010) && ({row_reg, col_reg}<19'b0110000110110010101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0110000110110010101)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0110000110110010110)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0110000110110010111) && ({row_reg, col_reg}<19'b0110000111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110000111001010001) && ({row_reg, col_reg}<19'b0110000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110000111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110000111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110001000000000000) && ({row_reg, col_reg}<19'b0110001000011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000011110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000011110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001000011110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110001000011110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001000011110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110001000011110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000011111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001000011111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001000011111011) && ({row_reg, col_reg}<19'b0110001000011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001000011111110) && ({row_reg, col_reg}<19'b0110001000100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000100000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001000100000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110001000100001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0110001000100001001) && ({row_reg, col_reg}<19'b0110001000100001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110001000100001011) && ({row_reg, col_reg}<19'b0110001000100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000100001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001000100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001000100010000) && ({row_reg, col_reg}<19'b0110001000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001000100011001) && ({row_reg, col_reg}<19'b0110001000100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000100011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0110001000100011100) && ({row_reg, col_reg}<19'b0110001000100011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001000100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000100100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110001000100100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110001000100100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110001000100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001000100100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110001000100100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110001000100100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110001000100100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0110001000100101000) && ({row_reg, col_reg}<19'b0110001000100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000100101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001000100101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110001000100101100) && ({row_reg, col_reg}<19'b0110001000100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001000100101111) && ({row_reg, col_reg}<19'b0110001000100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000100111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001000100111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001000100111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000100111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001000100111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001000100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000100111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0110001000101000000) && ({row_reg, col_reg}<19'b0110001000101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000101010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001000101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001000101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000101010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110001000101010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001000101010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000101010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110001000101011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110001000101011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001000101011010) && ({row_reg, col_reg}<19'b0110001000101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001000101011100) && ({row_reg, col_reg}<19'b0110001000101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001000101011110) && ({row_reg, col_reg}<19'b0110001000101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000101100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110001000101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001000101100010) && ({row_reg, col_reg}<19'b0110001000101100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110001000101100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001000101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001000101101000) && ({row_reg, col_reg}<19'b0110001000110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001000110001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001000110001111)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==19'b0110001000110010000)) color_data = 12'b011101111001;
		if(({row_reg, col_reg}==19'b0110001000110010001)) color_data = 12'b010000110110;
		if(({row_reg, col_reg}>=19'b0110001000110010010) && ({row_reg, col_reg}<19'b0110001000110010101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0110001000110010101)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0110001000110010110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110001000110010111) && ({row_reg, col_reg}<19'b0110001001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001001001010001) && ({row_reg, col_reg}<19'b0110001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110001001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110001001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110001010000000000) && ({row_reg, col_reg}<19'b0110001010011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010011110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110001010011110010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001010011110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010011110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110001010011110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001010011110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001010011110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110001010011111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001010011111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010011111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001010011111011) && ({row_reg, col_reg}<19'b0110001010011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001010011111101) && ({row_reg, col_reg}<19'b0110001010100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001010100001000) && ({row_reg, col_reg}<19'b0110001010100001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001010100001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001010100001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001010100001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001010100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001010100001110) && ({row_reg, col_reg}<19'b0110001010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010100011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110001010100011001) && ({row_reg, col_reg}<19'b0110001010100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001010100011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110001010100011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0110001010100011110) && ({row_reg, col_reg}<19'b0110001010100100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0110001010100100011) && ({row_reg, col_reg}<19'b0110001010100100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0110001010100100110) && ({row_reg, col_reg}<19'b0110001010100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010100101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001010100101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001010100101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0110001010100101011) && ({row_reg, col_reg}<19'b0110001010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010100101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001010100101111) && ({row_reg, col_reg}<19'b0110001010100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010100111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001010100111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010100111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010100111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001010100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010100111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0110001010101000000) && ({row_reg, col_reg}<19'b0110001010101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010101010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001010101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001010101010011) && ({row_reg, col_reg}<19'b0110001010101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010101010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110001010101010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010101011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001010101011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001010101011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110001010101011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001010101011100) && ({row_reg, col_reg}<19'b0110001010101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010101011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001010101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001010101100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0110001010101100001) && ({row_reg, col_reg}<19'b0110001010101100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010101100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001010101100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001010101100101) && ({row_reg, col_reg}<19'b0110001010110001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001010110001100) && ({row_reg, col_reg}<19'b0110001010110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001010110001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001010110001111)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==19'b0110001010110010000)) color_data = 12'b011001011000;
		if(({row_reg, col_reg}==19'b0110001010110010001)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==19'b0110001010110010010)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}>=19'b0110001010110010011) && ({row_reg, col_reg}<19'b0110001010110010101)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0110001010110010101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0110001010110010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110001010110010111) && ({row_reg, col_reg}<19'b0110001011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001011001010001) && ({row_reg, col_reg}<19'b0110001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110001011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110001011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110001100000000000) && ({row_reg, col_reg}<19'b0110001100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001100011110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110001100011110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110001100011110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100011110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0110001100011110100) && ({row_reg, col_reg}<19'b0110001100011110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001100011110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110001100011111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110001100011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001100011111011) && ({row_reg, col_reg}<19'b0110001100011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001100011111101) && ({row_reg, col_reg}<19'b0110001100100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001100100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001100100000100) && ({row_reg, col_reg}<19'b0110001100100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001100100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001100100001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001100100001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110001100100001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110001100100001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110001100100001100) && ({row_reg, col_reg}<19'b0110001100100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001100100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001100100011001) && ({row_reg, col_reg}<19'b0110001100100011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001100100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001100100011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0110001100100100000) && ({row_reg, col_reg}<19'b0110001100100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001100100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110001100100101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001100100101010) && ({row_reg, col_reg}<19'b0110001100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001100100111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110001100100111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001100100111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001100100111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001100100111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0110001100100111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001100100111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0110001100101000000) && ({row_reg, col_reg}<19'b0110001100101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001100101010001) && ({row_reg, col_reg}<19'b0110001100101010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001100101010011) && ({row_reg, col_reg}<19'b0110001100101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001100101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001100101010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100101010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0110001100101011000) && ({row_reg, col_reg}<19'b0110001100101011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001100101011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001100101011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001100101011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100101011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110001100101011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001100101011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001100101100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001100101100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110001100101100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001100101100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0110001100101100100) && ({row_reg, col_reg}<19'b0110001100110001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001100110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001100110001100) && ({row_reg, col_reg}<19'b0110001100110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001100110001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110001100110010000)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==19'b0110001100110010001)) color_data = 12'b000100010011;
		if(({row_reg, col_reg}==19'b0110001100110010010)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}==19'b0110001100110010011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0110001100110010100) && ({row_reg, col_reg}<19'b0110001100110010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110001100110010110) && ({row_reg, col_reg}<19'b0110001101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001101001010001) && ({row_reg, col_reg}<19'b0110001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110001101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110001101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110001110000000000) && ({row_reg, col_reg}<19'b0110001110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110011110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001110011110001) && ({row_reg, col_reg}<19'b0110001110011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110011110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110001110011110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001110011110101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001110011110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001110011110111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110001110011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001110011111001) && ({row_reg, col_reg}<19'b0110001110011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001110100000000) && ({row_reg, col_reg}<19'b0110001110100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001110100000011) && ({row_reg, col_reg}<19'b0110001110100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001110100000101) && ({row_reg, col_reg}<19'b0110001110100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001110100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001110100001001) && ({row_reg, col_reg}<19'b0110001110100001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110001110100001011) && ({row_reg, col_reg}<19'b0110001110100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001110100001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110001110100001111) && ({row_reg, col_reg}<19'b0110001110100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110100011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001110100011001) && ({row_reg, col_reg}<19'b0110001110100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110100011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001110100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001110100011101) && ({row_reg, col_reg}<19'b0110001110100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110100100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001110100100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110001110100100010) && ({row_reg, col_reg}<19'b0110001110100100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110001110100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001110100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001110100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001110100101001) && ({row_reg, col_reg}<19'b0110001110100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001110100101011) && ({row_reg, col_reg}<19'b0110001110100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001110100101101) && ({row_reg, col_reg}<19'b0110001110100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0110001110100111011) && ({row_reg, col_reg}<19'b0110001110100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001110100111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0110001110100111111) && ({row_reg, col_reg}<19'b0110001110101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110101010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110001110101010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001110101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001110101010101) && ({row_reg, col_reg}<19'b0110001110101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110101010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110001110101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001110101011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0110001110101011010) && ({row_reg, col_reg}<19'b0110001110101011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001110101011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0110001110101011110) && ({row_reg, col_reg}<19'b0110001110101100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001110101100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001110101100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110001110101100010) && ({row_reg, col_reg}<19'b0110001110110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001110110001001) && ({row_reg, col_reg}<19'b0110001110110001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110110001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001110110001100) && ({row_reg, col_reg}<19'b0110001110110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110110001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110001110110010000) && ({row_reg, col_reg}<19'b0110001110110010010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110001110110010010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0110001110110010011) && ({row_reg, col_reg}<19'b0110001110110010101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110001110110010101) && ({row_reg, col_reg}<19'b0110001110110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110001110110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110001110110011000) && ({row_reg, col_reg}<19'b0110001111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110001111001010001) && ({row_reg, col_reg}<19'b0110001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110001111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110001111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110010000000000000) && ({row_reg, col_reg}<19'b0110010000010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010000010101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110010000010101001) && ({row_reg, col_reg}<19'b0110010000010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010000010101011) && ({row_reg, col_reg}<19'b0110010000010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010000010101101) && ({row_reg, col_reg}<19'b0110010000010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010000010101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010000010110000) && ({row_reg, col_reg}<19'b0110010000010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010000010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010000010111001) && ({row_reg, col_reg}<19'b0110010000010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010000010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010000010111100) && ({row_reg, col_reg}<19'b0110010000011010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010000011010110) && ({row_reg, col_reg}<19'b0110010000011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010000011011000) && ({row_reg, col_reg}<19'b0110010000100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010000100111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110010000100111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110010000100111011) && ({row_reg, col_reg}<19'b0110010000100111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110010000100111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110010000100111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010000100111111) && ({row_reg, col_reg}<19'b0110010000101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010000101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110010000101011001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110010000101011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010000101011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0110010000101011100) && ({row_reg, col_reg}<19'b0110010000101011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110010000101011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110010000101011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0110010000101100000) && ({row_reg, col_reg}<19'b0110010000110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010000110010000) && ({row_reg, col_reg}<19'b0110010000110010100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110010000110010100) && ({row_reg, col_reg}<19'b0110010000110110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010000110110101) && ({row_reg, col_reg}<19'b0110010000110110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110010000110110111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110010000110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010000110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110010000110111010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0110010000110111011) && ({row_reg, col_reg}<19'b0110010000110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010000110111101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110010000110111110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0110010000110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0110010000111000000) && ({row_reg, col_reg}<19'b0110010001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010001001010001) && ({row_reg, col_reg}<19'b0110010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110010001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110010001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110010010000000000) && ({row_reg, col_reg}<19'b0110010010010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010010010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010010010101001) && ({row_reg, col_reg}<19'b0110010010010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010010010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110010010010101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110010010010101101) && ({row_reg, col_reg}<19'b0110010010010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010010010101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110010010010110000) && ({row_reg, col_reg}<19'b0110010010010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010010010110101) && ({row_reg, col_reg}<19'b0110010010010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010010010111001) && ({row_reg, col_reg}<19'b0110010010010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010010010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010010010111100) && ({row_reg, col_reg}<19'b0110010010010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010010010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010010011000000) && ({row_reg, col_reg}<19'b0110010010100111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010010100111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010010100111011) && ({row_reg, col_reg}<19'b0110010010100111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110010010100111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010010100111110) && ({row_reg, col_reg}<19'b0110010010101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010010101011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110010010101011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110010010101011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110010010101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110010010101011110) && ({row_reg, col_reg}<19'b0110010010101100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010010101100000) && ({row_reg, col_reg}<19'b0110010010110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010010110110000) && ({row_reg, col_reg}<19'b0110010010110111001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110010010110111001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==19'b0110010010110111010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=19'b0110010010110111011) && ({row_reg, col_reg}<19'b0110010010110111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110010010110111101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110010010110111110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0110010010110111111)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0110010010111000000) && ({row_reg, col_reg}<19'b0110010011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010011001010001) && ({row_reg, col_reg}<19'b0110010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110010011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110010011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110010100000000000) && ({row_reg, col_reg}<19'b0110010100010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010100010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010100010101001) && ({row_reg, col_reg}<19'b0110010100010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010100010101111) && ({row_reg, col_reg}<19'b0110010100010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010100010110010) && ({row_reg, col_reg}<19'b0110010100010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010100010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010100010111001) && ({row_reg, col_reg}<19'b0110010100010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010100010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110010100011000000) && ({row_reg, col_reg}<19'b0110010100101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010100101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010100101011001) && ({row_reg, col_reg}<19'b0110010100110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010100110110000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110010100110110001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110010100110110010) && ({row_reg, col_reg}<19'b0110010100110111000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110010100110111000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=19'b0110010100110111001) && ({row_reg, col_reg}<19'b0110010100110111011)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==19'b0110010100110111011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110010100110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110010100110111101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110010100110111110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==19'b0110010100110111111)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0110010100111000000) && ({row_reg, col_reg}<19'b0110010101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010101001010001) && ({row_reg, col_reg}<19'b0110010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110010101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110010101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110010110000000000) && ({row_reg, col_reg}<19'b0110010110010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010110010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010110010101001) && ({row_reg, col_reg}<19'b0110010110010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010110010110001) && ({row_reg, col_reg}<19'b0110010110010110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010110010110100) && ({row_reg, col_reg}<19'b0110010110010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010110010110110) && ({row_reg, col_reg}<19'b0110010110010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110010110010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110010110010111001) && ({row_reg, col_reg}<19'b0110010110010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010110010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010110011000000) && ({row_reg, col_reg}<19'b0110010110101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010110101011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110010110101011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010110101011010) && ({row_reg, col_reg}<19'b0110010110101011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110010110101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110010110101011110) && ({row_reg, col_reg}<19'b0110010110101100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110010110101100000) && ({row_reg, col_reg}<19'b0110010110110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010110110110000) && ({row_reg, col_reg}<19'b0110010110110110010)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110010110110110010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110010110110110011) && ({row_reg, col_reg}<19'b0110010110110110111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110010110110110111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110010110110111000)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==19'b0110010110110111001)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==19'b0110010110110111010)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==19'b0110010110110111011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0110010110110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110010110110111101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110010110110111110)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0110010110110111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110010110111000000) && ({row_reg, col_reg}<19'b0110010111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110010111001010001) && ({row_reg, col_reg}<19'b0110010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110010111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110010111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110011000000000000) && ({row_reg, col_reg}<19'b0110011000010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011000010101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011000010101110) && ({row_reg, col_reg}<19'b0110011000010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0110011000010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011000010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110011000010110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110011000010110011) && ({row_reg, col_reg}<19'b0110011000010110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011000010110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011000010110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011000010110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011000010111000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110011000010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011000010111010) && ({row_reg, col_reg}<19'b0110011000011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011000011011000) && ({row_reg, col_reg}<19'b0110011000011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011000011011010) && ({row_reg, col_reg}<19'b0110011000101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011000101011100) && ({row_reg, col_reg}<19'b0110011000101100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011000101100000) && ({row_reg, col_reg}<19'b0110011000110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011000110110000) && ({row_reg, col_reg}<19'b0110011000110110010)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0110011000110110010) && ({row_reg, col_reg}<19'b0110011000110110111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110011000110110111)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110011000110111000)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==19'b0110011000110111001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==19'b0110011000110111010)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==19'b0110011000110111011)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==19'b0110011000110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110011000110111101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110011000110111110)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0110011000110111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110011000111000000) && ({row_reg, col_reg}<19'b0110011001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011001001010001) && ({row_reg, col_reg}<19'b0110011001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110011001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110011001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110011010000000000) && ({row_reg, col_reg}<19'b0110011010010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011010010101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110011010010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0110011010010101110) && ({row_reg, col_reg}<19'b0110011010010110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011010010110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011010010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0110011010010110010) && ({row_reg, col_reg}<19'b0110011010010110100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011010010110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011010010110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011010010110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011010010110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011010010111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110011010010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110011010010111010) && ({row_reg, col_reg}<19'b0110011010011010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011010011010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011010011010110) && ({row_reg, col_reg}<19'b0110011010011011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110011010011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011010011011010) && ({row_reg, col_reg}<19'b0110011010100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011010100111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011010100111001) && ({row_reg, col_reg}<19'b0110011010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011010100111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011010101000000) && ({row_reg, col_reg}<19'b0110011010101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011010101011011) && ({row_reg, col_reg}<19'b0110011010101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011010101011101) && ({row_reg, col_reg}<19'b0110011010110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011010110110000) && ({row_reg, col_reg}<19'b0110011010110110101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110011010110110101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110011010110110110)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0110011010110110111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0110011010110111000)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==19'b0110011010110111001)) color_data = 12'b100101100111;
		if(({row_reg, col_reg}==19'b0110011010110111010)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==19'b0110011010110111011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0110011010110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110011010110111101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110011010110111110)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0110011010110111111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110011010111000000) && ({row_reg, col_reg}<19'b0110011011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011011001010001) && ({row_reg, col_reg}<19'b0110011011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110011011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110011011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110011100000000000) && ({row_reg, col_reg}<19'b0110011100010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011100010101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110011100010101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0110011100010101110) && ({row_reg, col_reg}<19'b0110011100010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011100010110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011100010110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011100010110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011100010110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110011100010110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110011100010110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011100010110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011100010111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110011100010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110011100010111010) && ({row_reg, col_reg}<19'b0110011100010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011100010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011100010111101) && ({row_reg, col_reg}<19'b0110011100011010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011100011010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110011100011010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110011100011010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110011100011011000) && ({row_reg, col_reg}<19'b0110011100011011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110011100011011010) && ({row_reg, col_reg}<19'b0110011100101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011100101011000) && ({row_reg, col_reg}<19'b0110011100101011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011100101011101) && ({row_reg, col_reg}<19'b0110011100110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011100110110000) && ({row_reg, col_reg}<19'b0110011100110110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110011100110110010) && ({row_reg, col_reg}<19'b0110011100110110100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110011100110110100)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110011100110110101)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0110011100110110110)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==19'b0110011100110110111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==19'b0110011100110111000)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==19'b0110011100110111001)) color_data = 12'b100101100111;
		if(({row_reg, col_reg}==19'b0110011100110111010)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==19'b0110011100110111011)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0110011100110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110011100110111101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110011100110111110)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==19'b0110011100110111111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110011100111000000) && ({row_reg, col_reg}<19'b0110011101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011101001010001) && ({row_reg, col_reg}<19'b0110011101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110011101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110011101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110011110000000000) && ({row_reg, col_reg}<19'b0110011110010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011110010101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110011110010101010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110011110010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011110010101100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110011110010101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110011110010101110)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==19'b0110011110010101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==19'b0110011110010110000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110011110010110001) && ({row_reg, col_reg}<19'b0110011110010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011110010110011) && ({row_reg, col_reg}<19'b0110011110010110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011110010110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110011110010110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011110010110111)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0110011110010111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110011110010111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011110010111010) && ({row_reg, col_reg}<19'b0110011110010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011110010111100) && ({row_reg, col_reg}<19'b0110011110010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110011110010111110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110011110010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011110011000000) && ({row_reg, col_reg}<19'b0110011110011010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011110011010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110011110011010101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==19'b0110011110011010110)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==19'b0110011110011010111)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==19'b0110011110011011000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==19'b0110011110011011001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==19'b0110011110011011010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110011110011011011) && ({row_reg, col_reg}<19'b0110011110101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110011110101011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110011110101011001) && ({row_reg, col_reg}<19'b0110011110110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011110110110000) && ({row_reg, col_reg}<19'b0110011110110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110011110110110011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110011110110110100)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0110011110110110101)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==19'b0110011110110110110)) color_data = 12'b011000010010;
		if(({row_reg, col_reg}==19'b0110011110110110111)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}==19'b0110011110110111000)) color_data = 12'b100101000101;
		if(({row_reg, col_reg}==19'b0110011110110111001)) color_data = 12'b101001010110;
		if(({row_reg, col_reg}==19'b0110011110110111010)) color_data = 12'b100001000100;
		if(({row_reg, col_reg}==19'b0110011110110111011)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}>=19'b0110011110110111100) && ({row_reg, col_reg}<19'b0110011110110111111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110011110110111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110011110111000000) && ({row_reg, col_reg}<19'b0110011111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110011111001010001) && ({row_reg, col_reg}<19'b0110011111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110011111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110011111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110100000000000000) && ({row_reg, col_reg}<19'b0110100000010100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100000010100100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100000010100101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100000010100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110100000010100111) && ({row_reg, col_reg}<19'b0110100000010101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100000010101001)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==19'b0110100000010101010)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0110100000010101011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110100000010101100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==19'b0110100000010101101)) color_data = 12'b110110101100;
		if(({row_reg, col_reg}==19'b0110100000010101110)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==19'b0110100000010101111)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=19'b0110100000010110000) && ({row_reg, col_reg}<19'b0110100000010110011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100000010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100000010110100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100000010110101)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==19'b0110100000010110110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==19'b0110100000010110111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=19'b0110100000010111000) && ({row_reg, col_reg}<19'b0110100000010111010)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0110100000010111010)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0110100000010111011) && ({row_reg, col_reg}<19'b0110100000010111101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110100000010111101) && ({row_reg, col_reg}<19'b0110100000011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100000011010000)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110100000011010001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100000011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100000011010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110100000011010100)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0110100000011010101)) color_data = 12'b011000010001;
		if(({row_reg, col_reg}==19'b0110100000011010110)) color_data = 12'b100100110011;
		if(({row_reg, col_reg}==19'b0110100000011010111)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==19'b0110100000011011000)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==19'b0110100000011011001)) color_data = 12'b011100010001;
		if(({row_reg, col_reg}==19'b0110100000011011010)) color_data = 12'b010100000000;
		if(({row_reg, col_reg}==19'b0110100000011011011)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0110100000011011100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==19'b0110100000011011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0110100000011011110) && ({row_reg, col_reg}<19'b0110100000011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100000011111000) && ({row_reg, col_reg}<19'b0110100000100000000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110100000100000000) && ({row_reg, col_reg}<19'b0110100000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100000100010001) && ({row_reg, col_reg}<19'b0110100000100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100000100011111) && ({row_reg, col_reg}<19'b0110100000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100000100101000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110100000100101001) && ({row_reg, col_reg}<19'b0110100000100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100000100110000) && ({row_reg, col_reg}<19'b0110100000100110010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110100000100110010) && ({row_reg, col_reg}<19'b0110100000100110100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110100000100110100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110100000100110101) && ({row_reg, col_reg}<19'b0110100000101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100000101000001) && ({row_reg, col_reg}<19'b0110100000101001111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100000101010000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110100000101010001) && ({row_reg, col_reg}<19'b0110100000101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100000101010111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100000101011000) && ({row_reg, col_reg}<19'b0110100000110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100000110110000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0110100000110110001) && ({row_reg, col_reg}<19'b0110100000110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110100000110110011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110100000110110100)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==19'b0110100000110110101)) color_data = 12'b011100000001;
		if(({row_reg, col_reg}==19'b0110100000110110110)) color_data = 12'b101100100011;
		if(({row_reg, col_reg}>=19'b0110100000110110111) && ({row_reg, col_reg}<19'b0110100000110111001)) color_data = 12'b110001000101;
		if(({row_reg, col_reg}==19'b0110100000110111001)) color_data = 12'b110000110100;
		if(({row_reg, col_reg}==19'b0110100000110111010)) color_data = 12'b100100100011;
		if(({row_reg, col_reg}==19'b0110100000110111011)) color_data = 12'b011000010000;
		if(({row_reg, col_reg}==19'b0110100000110111100)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}>=19'b0110100000110111101) && ({row_reg, col_reg}<19'b0110100000110111111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110100000110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0110100000111000000) && ({row_reg, col_reg}<19'b0110100001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100001001010001) && ({row_reg, col_reg}<19'b0110100001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110100001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110100010000000000) && ({row_reg, col_reg}<19'b0110100010010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100010010100001) && ({row_reg, col_reg}<19'b0110100010010101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100010010101001)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0110100010010101010)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0110100010010101011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100010010101100)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==19'b0110100010010101101)) color_data = 12'b101110001011;
		if(({row_reg, col_reg}==19'b0110100010010101110)) color_data = 12'b101101111010;
		if(({row_reg, col_reg}==19'b0110100010010101111)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0110100010010110000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0110100010010110001) && ({row_reg, col_reg}<19'b0110100010010110011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100010010110011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100010010110100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100010010110101)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0110100010010110110)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==19'b0110100010010110111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=19'b0110100010010111000) && ({row_reg, col_reg}<19'b0110100010010111010)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0110100010010111010)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0110100010010111011) && ({row_reg, col_reg}<19'b0110100010010111101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110100010010111101) && ({row_reg, col_reg}<19'b0110100010010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110100010010111111) && ({row_reg, col_reg}<19'b0110100010011010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100010011010011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110100010011010100)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==19'b0110100010011010101)) color_data = 12'b100000100010;
		if(({row_reg, col_reg}==19'b0110100010011010110)) color_data = 12'b101100110010;
		if(({row_reg, col_reg}>=19'b0110100010011010111) && ({row_reg, col_reg}<19'b0110100010011011001)) color_data = 12'b110000110011;
		if(({row_reg, col_reg}==19'b0110100010011011001)) color_data = 12'b100100010001;
		if(({row_reg, col_reg}==19'b0110100010011011010)) color_data = 12'b010100000000;
		if(({row_reg, col_reg}==19'b0110100010011011011)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0110100010011011100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110100010011011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100010011011110) && ({row_reg, col_reg}<19'b0110100010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100010011111000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110100010011111001) && ({row_reg, col_reg}<19'b0110100010011111011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110100010011111011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110100010011111100) && ({row_reg, col_reg}<19'b0110100010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100010100010000) && ({row_reg, col_reg}<19'b0110100010100100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100010100100000) && ({row_reg, col_reg}<19'b0110100010100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100010100101100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110100010100101101) && ({row_reg, col_reg}<19'b0110100010100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110100010100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100010100110001) && ({row_reg, col_reg}<19'b0110100010100110011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110100010100110011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110100010100110100) && ({row_reg, col_reg}<19'b0110100010100110110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110100010100110110) && ({row_reg, col_reg}<19'b0110100010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100010101000000) && ({row_reg, col_reg}<19'b0110100010101010000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110100010101010000) && ({row_reg, col_reg}<19'b0110100010101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100010101010010) && ({row_reg, col_reg}<19'b0110100010101010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100010101010110) && ({row_reg, col_reg}<19'b0110100010110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100010110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110100010110110010)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==19'b0110100010110110011)) color_data = 12'b010100010000;
		if(({row_reg, col_reg}==19'b0110100010110110100)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==19'b0110100010110110101)) color_data = 12'b101000100010;
		if(({row_reg, col_reg}==19'b0110100010110110110)) color_data = 12'b110000100011;
		if(({row_reg, col_reg}==19'b0110100010110110111)) color_data = 12'b110100110011;
		if(({row_reg, col_reg}==19'b0110100010110111000)) color_data = 12'b110100100011;
		if(({row_reg, col_reg}==19'b0110100010110111001)) color_data = 12'b110100110100;
		if(({row_reg, col_reg}==19'b0110100010110111010)) color_data = 12'b110001000100;
		if(({row_reg, col_reg}==19'b0110100010110111011)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==19'b0110100010110111100)) color_data = 12'b011000100000;
		if(({row_reg, col_reg}==19'b0110100010110111101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110100010110111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100010110111111) && ({row_reg, col_reg}<19'b0110100011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100011001010001) && ({row_reg, col_reg}<19'b0110100011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110100011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110100100000000000) && ({row_reg, col_reg}<19'b0110100100010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100100010100001) && ({row_reg, col_reg}<19'b0110100100010100111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100100010100111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100100010101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110100100010101001) && ({row_reg, col_reg}<19'b0110100100010101011)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0110100100010101011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100100010101100)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==19'b0110100100010101101)) color_data = 12'b101110001010;
		if(({row_reg, col_reg}==19'b0110100100010101110)) color_data = 12'b101001101001;
		if(({row_reg, col_reg}==19'b0110100100010101111)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0110100100010110000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0110100100010110001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110100100010110010) && ({row_reg, col_reg}<19'b0110100100010110100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100100010110100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100100010110101)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==19'b0110100100010110110)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==19'b0110100100010110111)) color_data = 12'b110010111101;
		if(({row_reg, col_reg}==19'b0110100100010111000)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=19'b0110100100010111001) && ({row_reg, col_reg}<19'b0110100100010111011)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0110100100010111011) && ({row_reg, col_reg}<19'b0110100100010111101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110100100010111101) && ({row_reg, col_reg}<19'b0110100100010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110100100010111111) && ({row_reg, col_reg}<19'b0110100100011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100100011010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110100100011010011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==19'b0110100100011010100)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}==19'b0110100100011010101)) color_data = 12'b100100110011;
		if(({row_reg, col_reg}==19'b0110100100011010110)) color_data = 12'b101100110011;
		if(({row_reg, col_reg}==19'b0110100100011010111)) color_data = 12'b110000110011;
		if(({row_reg, col_reg}==19'b0110100100011011000)) color_data = 12'b110101000100;
		if(({row_reg, col_reg}==19'b0110100100011011001)) color_data = 12'b101000100010;
		if(({row_reg, col_reg}==19'b0110100100011011010)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==19'b0110100100011011011)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0110100100011011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110100100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100100011011110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100100011011111)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110100100011100000) && ({row_reg, col_reg}<19'b0110100100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100100011111000) && ({row_reg, col_reg}<19'b0110100100011111100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110100100011111100) && ({row_reg, col_reg}<19'b0110100100100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100100100010001) && ({row_reg, col_reg}<19'b0110100100100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100100100011111) && ({row_reg, col_reg}<19'b0110100100100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100100100101010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110100100100101011) && ({row_reg, col_reg}<19'b0110100100100110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110100100100110000) && ({row_reg, col_reg}<19'b0110100100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100100100110011) && ({row_reg, col_reg}<19'b0110100100100111000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110100100100111000) && ({row_reg, col_reg}<19'b0110100100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100100101000000) && ({row_reg, col_reg}<19'b0110100100101010000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110100100101010000) && ({row_reg, col_reg}<19'b0110100100101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100100101010010) && ({row_reg, col_reg}<19'b0110100100101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110100100101010110) && ({row_reg, col_reg}<19'b0110100100110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100100110110001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0110100100110110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==19'b0110100100110110011)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==19'b0110100100110110100)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==19'b0110100100110110101)) color_data = 12'b110001000100;
		if(({row_reg, col_reg}==19'b0110100100110110110)) color_data = 12'b110000110100;
		if(({row_reg, col_reg}>=19'b0110100100110110111) && ({row_reg, col_reg}<19'b0110100100110111001)) color_data = 12'b110000100011;
		if(({row_reg, col_reg}==19'b0110100100110111001)) color_data = 12'b110100110100;
		if(({row_reg, col_reg}==19'b0110100100110111010)) color_data = 12'b110101010101;
		if(({row_reg, col_reg}==19'b0110100100110111011)) color_data = 12'b110001010101;
		if(({row_reg, col_reg}==19'b0110100100110111100)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==19'b0110100100110111101)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==19'b0110100100110111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100100110111111) && ({row_reg, col_reg}<19'b0110100101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100101001010001) && ({row_reg, col_reg}<19'b0110100101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110100101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110100110000000000) && ({row_reg, col_reg}<19'b0110100110010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100110010100001) && ({row_reg, col_reg}<19'b0110100110010100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100110010100110)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0110100110010100111)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0110100110010101000)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}>=19'b0110100110010101001) && ({row_reg, col_reg}<19'b0110100110010101011)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==19'b0110100110010101011)) color_data = 12'b011000110101;
		if(({row_reg, col_reg}==19'b0110100110010101100)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==19'b0110100110010101101)) color_data = 12'b110110101100;
		if(({row_reg, col_reg}==19'b0110100110010101110)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==19'b0110100110010101111)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0110100110010110000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110100110010110001) && ({row_reg, col_reg}<19'b0110100110010110100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100110010110100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100110010110101)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==19'b0110100110010110110)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==19'b0110100110010110111)) color_data = 12'b110110111101;
		if(({row_reg, col_reg}>=19'b0110100110010111000) && ({row_reg, col_reg}<19'b0110100110010111010)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0110100110010111010)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0110100110010111011) && ({row_reg, col_reg}<19'b0110100110010111110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110100110010111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110100110010111111) && ({row_reg, col_reg}<19'b0110100110011010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100110011010001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100110011010010)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==19'b0110100110011010011)) color_data = 12'b011101000100;
		if(({row_reg, col_reg}==19'b0110100110011010100)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==19'b0110100110011010101)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}>=19'b0110100110011010110) && ({row_reg, col_reg}<19'b0110100110011011000)) color_data = 12'b101100110011;
		if(({row_reg, col_reg}==19'b0110100110011011000)) color_data = 12'b110001000100;
		if(({row_reg, col_reg}==19'b0110100110011011001)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==19'b0110100110011011010)) color_data = 12'b011100010001;
		if(({row_reg, col_reg}==19'b0110100110011011011)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==19'b0110100110011011100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110100110011011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100110011011110) && ({row_reg, col_reg}<19'b0110100110011100000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110100110011100000) && ({row_reg, col_reg}<19'b0110100110011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100110011111011) && ({row_reg, col_reg}<19'b0110100110011111101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110100110011111101) && ({row_reg, col_reg}<19'b0110100110100000000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110100110100000000) && ({row_reg, col_reg}<19'b0110100110100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100110100010001) && ({row_reg, col_reg}<19'b0110100110100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100110100011111) && ({row_reg, col_reg}<19'b0110100110100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100110100101010) && ({row_reg, col_reg}<19'b0110100110100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110100110100101101) && ({row_reg, col_reg}<19'b0110100110100110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100110100110101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110100110100110110) && ({row_reg, col_reg}<19'b0110100110100111000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110100110100111000) && ({row_reg, col_reg}<19'b0110100110101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100110101000000) && ({row_reg, col_reg}<19'b0110100110101001111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110100110101001111) && ({row_reg, col_reg}<19'b0110100110110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110100110110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110100110110110010)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==19'b0110100110110110011)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==19'b0110100110110110100)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==19'b0110100110110110101)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}==19'b0110100110110110110)) color_data = 12'b101100110011;
		if(({row_reg, col_reg}>=19'b0110100110110110111) && ({row_reg, col_reg}<19'b0110100110110111001)) color_data = 12'b101100100011;
		if(({row_reg, col_reg}==19'b0110100110110111001)) color_data = 12'b110001000100;
		if(({row_reg, col_reg}==19'b0110100110110111010)) color_data = 12'b110001010101;
		if(({row_reg, col_reg}==19'b0110100110110111011)) color_data = 12'b101101010101;
		if(({row_reg, col_reg}==19'b0110100110110111100)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==19'b0110100110110111101)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==19'b0110100110110111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110100110110111111) && ({row_reg, col_reg}<19'b0110100111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110100111001010001) && ({row_reg, col_reg}<19'b0110100111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110100111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110100111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110101000000000000) && ({row_reg, col_reg}<19'b0110101000010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101000010100001) && ({row_reg, col_reg}<19'b0110101000010100110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101000010100110)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==19'b0110101000010100111)) color_data = 12'b010101000110;
		if(({row_reg, col_reg}==19'b0110101000010101000)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}>=19'b0110101000010101001) && ({row_reg, col_reg}<19'b0110101000010101011)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0110101000010101011)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==19'b0110101000010101100)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}==19'b0110101000010101101)) color_data = 12'b110110101101;
		if(({row_reg, col_reg}==19'b0110101000010101110)) color_data = 12'b100101101001;
		if(({row_reg, col_reg}==19'b0110101000010101111)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0110101000010110000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110101000010110001) && ({row_reg, col_reg}<19'b0110101000010110011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101000010110011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110101000010110100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0110101000010110101)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==19'b0110101000010110110)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0110101000010110111)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==19'b0110101000010111000)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0110101000010111001) && ({row_reg, col_reg}<19'b0110101000010111111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110101000010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110101000011000000) && ({row_reg, col_reg}<19'b0110101000011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101000011010000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101000011010001)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==19'b0110101000011010010)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==19'b0110101000011010011)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==19'b0110101000011010100)) color_data = 12'b100101010101;
		if(({row_reg, col_reg}==19'b0110101000011010101)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}>=19'b0110101000011010110) && ({row_reg, col_reg}<19'b0110101000011011000)) color_data = 12'b101000110010;
		if(({row_reg, col_reg}>=19'b0110101000011011000) && ({row_reg, col_reg}<19'b0110101000011011010)) color_data = 12'b101101000011;
		if(({row_reg, col_reg}==19'b0110101000011011010)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==19'b0110101000011011011)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==19'b0110101000011011100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==19'b0110101000011011101)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=19'b0110101000011011110) && ({row_reg, col_reg}<19'b0110101000011100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110101000011100000) && ({row_reg, col_reg}<19'b0110101000011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101000011111011) && ({row_reg, col_reg}<19'b0110101000100000000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110101000100000000) && ({row_reg, col_reg}<19'b0110101000100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101000100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110101000100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110101000100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110101000100101100) && ({row_reg, col_reg}<19'b0110101000100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101000100110000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110101000100110001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110101000100110010) && ({row_reg, col_reg}<19'b0110101000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101000100110110) && ({row_reg, col_reg}<19'b0110101000100111000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110101000100111000) && ({row_reg, col_reg}<19'b0110101000101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101000101000001) && ({row_reg, col_reg}<19'b0110101000101001111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101000101010000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110101000101010001) && ({row_reg, col_reg}<19'b0110101000110110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101000110110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110101000110110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==19'b0110101000110110011)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==19'b0110101000110110100)) color_data = 12'b011000010001;
		if(({row_reg, col_reg}==19'b0110101000110110101)) color_data = 12'b100000100010;
		if(({row_reg, col_reg}==19'b0110101000110110110)) color_data = 12'b101000100010;
		if(({row_reg, col_reg}==19'b0110101000110110111)) color_data = 12'b101000100011;
		if(({row_reg, col_reg}==19'b0110101000110111000)) color_data = 12'b110000110100;
		if(({row_reg, col_reg}==19'b0110101000110111001)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}==19'b0110101000110111010)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==19'b0110101000110111011)) color_data = 12'b100000110010;
		if(({row_reg, col_reg}==19'b0110101000110111100)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==19'b0110101000110111101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110101000110111110) && ({row_reg, col_reg}<19'b0110101001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101001001010001) && ({row_reg, col_reg}<19'b0110101001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110101001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110101010000000000) && ({row_reg, col_reg}<19'b0110101010010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101010010100001) && ({row_reg, col_reg}<19'b0110101010010100101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101010010100101)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0110101010010100110)) color_data = 12'b010101000110;
		if(({row_reg, col_reg}==19'b0110101010010100111)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}==19'b0110101010010101000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==19'b0110101010010101001)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0110101010010101010)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}==19'b0110101010010101011)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}>=19'b0110101010010101100) && ({row_reg, col_reg}<19'b0110101010010101110)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0110101010010101110)) color_data = 12'b100001000111;
		if(({row_reg, col_reg}>=19'b0110101010010101111) && ({row_reg, col_reg}<19'b0110101010010110010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110101010010110010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0110101010010110011)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==19'b0110101010010110100)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==19'b0110101010010110101)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==19'b0110101010010110110)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0110101010010110111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=19'b0110101010010111000) && ({row_reg, col_reg}<19'b0110101010011000000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110101010011000000) && ({row_reg, col_reg}<19'b0110101010011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101010011010000)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0110101010011010001)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==19'b0110101010011010010)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==19'b0110101010011010011)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==19'b0110101010011010100)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}==19'b0110101010011010101)) color_data = 12'b011100100010;
		if(({row_reg, col_reg}==19'b0110101010011010110)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==19'b0110101010011010111)) color_data = 12'b101001000011;
		if(({row_reg, col_reg}==19'b0110101010011011000)) color_data = 12'b101000110011;
		if(({row_reg, col_reg}==19'b0110101010011011001)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}==19'b0110101010011011010)) color_data = 12'b101001100101;
		if(({row_reg, col_reg}==19'b0110101010011011011)) color_data = 12'b100101010101;
		if(({row_reg, col_reg}==19'b0110101010011011100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==19'b0110101010011011101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0110101010011011110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110101010011011111) && ({row_reg, col_reg}<19'b0110101010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101010011111000) && ({row_reg, col_reg}<19'b0110101010011111010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110101010011111010) && ({row_reg, col_reg}<19'b0110101010011111100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110101010011111100) && ({row_reg, col_reg}<19'b0110101010100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101010100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110101010100101010)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110101010100101011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0110101010100101100) && ({row_reg, col_reg}<19'b0110101010100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101010100101110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110101010100101111)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0110101010100110000)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110101010100110001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110101010100110010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110101010100110011) && ({row_reg, col_reg}<19'b0110101010100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101010100110111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110101010100111000) && ({row_reg, col_reg}<19'b0110101010101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101010101010000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110101010101010001) && ({row_reg, col_reg}<19'b0110101010110110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101010110110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110101010110110011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110101010110110100)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0110101010110110101)) color_data = 12'b010100000000;
		if(({row_reg, col_reg}==19'b0110101010110110110)) color_data = 12'b011100000001;
		if(({row_reg, col_reg}==19'b0110101010110110111)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==19'b0110101010110111000)) color_data = 12'b101101000101;
		if(({row_reg, col_reg}==19'b0110101010110111001)) color_data = 12'b101101000100;
		if(({row_reg, col_reg}==19'b0110101010110111010)) color_data = 12'b100000110011;
		if(({row_reg, col_reg}==19'b0110101010110111011)) color_data = 12'b010100010000;
		if(({row_reg, col_reg}==19'b0110101010110111100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110101010110111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110101010110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101010110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0110101010111000000) && ({row_reg, col_reg}<19'b0110101011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101011001010001) && ({row_reg, col_reg}<19'b0110101011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110101011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110101100000000000) && ({row_reg, col_reg}<19'b0110101100010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101100010100001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101100010100010)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0110101100010100011) && ({row_reg, col_reg}<19'b0110101100010100101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101100010100101)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==19'b0110101100010100110)) color_data = 12'b011101101000;
		if(({row_reg, col_reg}==19'b0110101100010100111)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}>=19'b0110101100010101000) && ({row_reg, col_reg}<19'b0110101100010101011)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0110101100010101011)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0110101100010101100)) color_data = 12'b110110101100;
		if(({row_reg, col_reg}==19'b0110101100010101101)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}==19'b0110101100010101110)) color_data = 12'b011101000110;
		if(({row_reg, col_reg}>=19'b0110101100010101111) && ({row_reg, col_reg}<19'b0110101100010110001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110101100010110001)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==19'b0110101100010110010)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==19'b0110101100010110011)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==19'b0110101100010110100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==19'b0110101100010110101)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}>=19'b0110101100010110110) && ({row_reg, col_reg}<19'b0110101100010111000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=19'b0110101100010111000) && ({row_reg, col_reg}<19'b0110101100011000000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110101100011000000) && ({row_reg, col_reg}<19'b0110101100011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101100011010000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101100011010001)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==19'b0110101100011010010)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==19'b0110101100011010011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==19'b0110101100011010100)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==19'b0110101100011010101)) color_data = 12'b010100010000;
		if(({row_reg, col_reg}==19'b0110101100011010110)) color_data = 12'b100000110010;
		if(({row_reg, col_reg}==19'b0110101100011010111)) color_data = 12'b101101010100;
		if(({row_reg, col_reg}==19'b0110101100011011000)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}==19'b0110101100011011001)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}==19'b0110101100011011010)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}==19'b0110101100011011011)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==19'b0110101100011011100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==19'b0110101100011011101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110101100011011110) && ({row_reg, col_reg}<19'b0110101100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101100011111000) && ({row_reg, col_reg}<19'b0110101100011111010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110101100011111010) && ({row_reg, col_reg}<19'b0110101100011111100)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110101100011111100)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}>=19'b0110101100011111101) && ({row_reg, col_reg}<19'b0110101100011111111)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0110101100011111111)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}>=19'b0110101100100000000) && ({row_reg, col_reg}<19'b0110101100100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101100100101001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110101100100101010)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110101100100101011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110101100100101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101100100101101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0110101100100101110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==19'b0110101100100101111)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==19'b0110101100100110000)) color_data = 12'b001000110011;
		if(({row_reg, col_reg}==19'b0110101100100110001)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110101100100110010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110101100100110011) && ({row_reg, col_reg}<19'b0110101100101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101100101010001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110101100101010010)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0110101100101010011) && ({row_reg, col_reg}<19'b0110101100101010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110101100101010101)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110101100101010110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110101100101010111) && ({row_reg, col_reg}<19'b0110101100110110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101100110110010) && ({row_reg, col_reg}<19'b0110101100110110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110101100110110100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110101100110110101)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0110101100110110110)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==19'b0110101100110110111)) color_data = 12'b010100000000;
		if(({row_reg, col_reg}==19'b0110101100110111000)) color_data = 12'b101101000101;
		if(({row_reg, col_reg}==19'b0110101100110111001)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==19'b0110101100110111010)) color_data = 12'b100000110011;
		if(({row_reg, col_reg}==19'b0110101100110111011)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}>=19'b0110101100110111100) && ({row_reg, col_reg}<19'b0110101100110111110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110101100110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101100110111111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0110101100111000000) && ({row_reg, col_reg}<19'b0110101101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101101001010001) && ({row_reg, col_reg}<19'b0110101101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110101101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110101110000000000) && ({row_reg, col_reg}<19'b0110101110010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101110010100001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101110010100010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0110101110010100011) && ({row_reg, col_reg}<19'b0110101110010100101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101110010100101)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==19'b0110101110010100110)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==19'b0110101110010100111)) color_data = 12'b110111001110;
		if(({row_reg, col_reg}>=19'b0110101110010101000) && ({row_reg, col_reg}<19'b0110101110010101010)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0110101110010101010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==19'b0110101110010101011)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0110101110010101100)) color_data = 12'b110110101100;
		if(({row_reg, col_reg}==19'b0110101110010101101)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}==19'b0110101110010101110)) color_data = 12'b011101000110;
		if(({row_reg, col_reg}==19'b0110101110010101111)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110101110010110000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110101110010110001)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0110101110010110010)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0110101110010110011)) color_data = 12'b110010111101;
		if(({row_reg, col_reg}==19'b0110101110010110100)) color_data = 12'b110111001101;
		if(({row_reg, col_reg}==19'b0110101110010110101)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0110101110010110110)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0110101110010110111)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}>=19'b0110101110010111000) && ({row_reg, col_reg}<19'b0110101110011000000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110101110011000000) && ({row_reg, col_reg}<19'b0110101110011010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101110011010001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110101110011010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0110101110011010011) && ({row_reg, col_reg}<19'b0110101110011010101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110101110011010101)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0110101110011010110)) color_data = 12'b011100110010;
		if(({row_reg, col_reg}==19'b0110101110011010111)) color_data = 12'b101101110101;
		if(({row_reg, col_reg}>=19'b0110101110011011000) && ({row_reg, col_reg}<19'b0110101110011011010)) color_data = 12'b100101010011;
		if(({row_reg, col_reg}==19'b0110101110011011010)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==19'b0110101110011011011)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==19'b0110101110011011100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110101110011011101) && ({row_reg, col_reg}<19'b0110101110011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101110011011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110101110011100000) && ({row_reg, col_reg}<19'b0110101110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101110011111001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110101110011111010)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110101110011111011)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110101110011111100)) color_data = 12'b001101100101;
		if(({row_reg, col_reg}==19'b0110101110011111101)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110101110011111110)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0110101110011111111)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}>=19'b0110101110100000000) && ({row_reg, col_reg}<19'b0110101110100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101110100101010)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}>=19'b0110101110100101011) && ({row_reg, col_reg}<19'b0110101110100101101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110101110100101101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0110101110100101110)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==19'b0110101110100101111)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==19'b0110101110100110000)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==19'b0110101110100110001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0110101110100110010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110101110100110011) && ({row_reg, col_reg}<19'b0110101110101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110101110101010001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110101110101010010)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}>=19'b0110101110101010011) && ({row_reg, col_reg}<19'b0110101110101010101)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==19'b0110101110101010101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==19'b0110101110101010110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110101110101010111) && ({row_reg, col_reg}<19'b0110101110110110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101110110110010) && ({row_reg, col_reg}<19'b0110101110110110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110101110110110100) && ({row_reg, col_reg}<19'b0110101110110110110)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110101110110110110) && ({row_reg, col_reg}<19'b0110101110110111000)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==19'b0110101110110111000)) color_data = 12'b100101000101;
		if(({row_reg, col_reg}==19'b0110101110110111001)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==19'b0110101110110111010)) color_data = 12'b011100110100;
		if(({row_reg, col_reg}==19'b0110101110110111011)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==19'b0110101110110111100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110101110110111101) && ({row_reg, col_reg}<19'b0110101111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110101111001010001) && ({row_reg, col_reg}<19'b0110101111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110101111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110101111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110110000000000000) && ({row_reg, col_reg}<19'b0110110000010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000010100000)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0110110000010100001) && ({row_reg, col_reg}<19'b0110110000010100101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110110000010100101)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==19'b0110110000010100110)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}==19'b0110110000010100111)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0110110000010101000)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0110110000010101001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==19'b0110110000010101010)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0110110000010101011)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0110110000010101100)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==19'b0110110000010101101)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0110110000010101110)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0110110000010101111)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110110000010110000)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0110110000010110001)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==19'b0110110000010110010)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}>=19'b0110110000010110011) && ({row_reg, col_reg}<19'b0110110000010110101)) color_data = 12'b111011001110;
		if(({row_reg, col_reg}==19'b0110110000010110101)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}==19'b0110110000010110110)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==19'b0110110000010110111)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=19'b0110110000010111000) && ({row_reg, col_reg}<19'b0110110000010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110110000010111111) && ({row_reg, col_reg}<19'b0110110000011010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000011010001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110110000011010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0110110000011010011) && ({row_reg, col_reg}<19'b0110110000011010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110000011010101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110110000011010110)) color_data = 12'b011000110001;
		if(({row_reg, col_reg}>=19'b0110110000011010111) && ({row_reg, col_reg}<19'b0110110000011011001)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}==19'b0110110000011011001)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==19'b0110110000011011010)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==19'b0110110000011011011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110110000011011100) && ({row_reg, col_reg}<19'b0110110000011011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110000011011110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110110000011011111) && ({row_reg, col_reg}<19'b0110110000011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110000011110001) && ({row_reg, col_reg}<19'b0110110000011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110000011110011) && ({row_reg, col_reg}<19'b0110110000011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000011110110)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==19'b0110110000011110111)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==19'b0110110000011111000)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==19'b0110110000011111001)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110110000011111010)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==19'b0110110000011111011)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}>=19'b0110110000011111100) && ({row_reg, col_reg}<19'b0110110000011111110)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==19'b0110110000011111110)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==19'b0110110000011111111)) color_data = 12'b110011111110;
		if(({row_reg, col_reg}==19'b0110110000100000000)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}>=19'b0110110000100000001) && ({row_reg, col_reg}<19'b0110110000100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000100000011)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110110000100000100)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}>=19'b0110110000100000101) && ({row_reg, col_reg}<19'b0110110000100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000100000111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110110000100001000) && ({row_reg, col_reg}<19'b0110110000100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000100001010)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110110000100001011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110110000100001100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110110000100001101)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}>=19'b0110110000100001110) && ({row_reg, col_reg}<19'b0110110000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110000100011000) && ({row_reg, col_reg}<19'b0110110000100011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110000100011100) && ({row_reg, col_reg}<19'b0110110000100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000100011110)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110110000100011111)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==19'b0110110000100100000)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110110000100100001)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110110000100100010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110000100100011)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0110110000100100100) && ({row_reg, col_reg}<19'b0110110000100100110)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0110110000100100110)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110110000100100111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110000100101000)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110110000100101001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110000100101010) && ({row_reg, col_reg}<19'b0110110000100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000100101101)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110110000100101110)) color_data = 12'b010101100101;
		if(({row_reg, col_reg}==19'b0110110000100101111)) color_data = 12'b100110111001;
		if(({row_reg, col_reg}==19'b0110110000100110000)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}>=19'b0110110000100110001) && ({row_reg, col_reg}<19'b0110110000100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000100110011)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110110000100110100) && ({row_reg, col_reg}<19'b0110110000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000100110110)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0110110000100110111) && ({row_reg, col_reg}<19'b0110110000100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000100111001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110110000100111010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110110000100111011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110110000100111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110000100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000100111110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110110000100111111) && ({row_reg, col_reg}<19'b0110110000101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110000101000100) && ({row_reg, col_reg}<19'b0110110000101000110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110110000101000110) && ({row_reg, col_reg}<19'b0110110000101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000101001010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110000101001011) && ({row_reg, col_reg}<19'b0110110000101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000101010010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110000101010011)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==19'b0110110000101010100)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==19'b0110110000101010101)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==19'b0110110000101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000101010111)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}>=19'b0110110000101011000) && ({row_reg, col_reg}<19'b0110110000101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110000101011100) && ({row_reg, col_reg}<19'b0110110000101011110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110000101011110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110000101011111) && ({row_reg, col_reg}<19'b0110110000101100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110000101100010) && ({row_reg, col_reg}<19'b0110110000101100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110000101100101) && ({row_reg, col_reg}<19'b0110110000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110000101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110000101111001) && ({row_reg, col_reg}<19'b0110110000110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110000110110011) && ({row_reg, col_reg}<19'b0110110000110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110110000110110101) && ({row_reg, col_reg}<19'b0110110000110111011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110110000110111011) && ({row_reg, col_reg}<19'b0110110000110111101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110110000110111101) && ({row_reg, col_reg}<19'b0110110001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110001001010001) && ({row_reg, col_reg}<19'b0110110001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110110001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110110001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110110010000000000) && ({row_reg, col_reg}<19'b0110110010010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010010100000)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0110110010010100001) && ({row_reg, col_reg}<19'b0110110010010100101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110110010010100101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0110110010010100110)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==19'b0110110010010100111)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}>=19'b0110110010010101000) && ({row_reg, col_reg}<19'b0110110010010101010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0110110010010101010)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0110110010010101011)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0110110010010101100) && ({row_reg, col_reg}<19'b0110110010010101111)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110110010010101111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110110010010110000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110110010010110001)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0110110010010110010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=19'b0110110010010110011) && ({row_reg, col_reg}<19'b0110110010010110101)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==19'b0110110010010110101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==19'b0110110010010110110)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0110110010010110111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110110010010111000) && ({row_reg, col_reg}<19'b0110110010010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110110010010111111) && ({row_reg, col_reg}<19'b0110110010011010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010011010001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110110010011010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=19'b0110110010011010011) && ({row_reg, col_reg}<19'b0110110010011010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110010011010101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==19'b0110110010011010110)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==19'b0110110010011010111)) color_data = 12'b100001100100;
		if(({row_reg, col_reg}==19'b0110110010011011000)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==19'b0110110010011011001)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==19'b0110110010011011010)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==19'b0110110010011011011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=19'b0110110010011011100) && ({row_reg, col_reg}<19'b0110110010011011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110010011011110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110110010011011111) && ({row_reg, col_reg}<19'b0110110010011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110010011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110010011110011) && ({row_reg, col_reg}<19'b0110110010011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010011110101)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110110010011110110)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==19'b0110110010011110111)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=19'b0110110010011111000) && ({row_reg, col_reg}<19'b0110110010011111011)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0110110010011111011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==19'b0110110010011111100)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}>=19'b0110110010011111101) && ({row_reg, col_reg}<19'b0110110010011111111)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==19'b0110110010011111111)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110110010100000000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110110010100000001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110010100000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110010100000011) && ({row_reg, col_reg}<19'b0110110010100000101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110010100000101) && ({row_reg, col_reg}<19'b0110110010100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010100001000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110010100001001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110010100001010)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}>=19'b0110110010100001011) && ({row_reg, col_reg}<19'b0110110010100001101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110110010100001101)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}>=19'b0110110010100001110) && ({row_reg, col_reg}<19'b0110110010100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110010100100000) && ({row_reg, col_reg}<19'b0110110010100101001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110010100101001) && ({row_reg, col_reg}<19'b0110110010100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010100101101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110010100101110)) color_data = 12'b010001100100;
		if(({row_reg, col_reg}==19'b0110110010100101111)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==19'b0110110010100110000)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}>=19'b0110110010100110001) && ({row_reg, col_reg}<19'b0110110010100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010100110011)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110110010100110100) && ({row_reg, col_reg}<19'b0110110010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010100110110)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0110110010100110111) && ({row_reg, col_reg}<19'b0110110010100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010100111001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110110010100111010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110110010100111011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110110010100111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110010100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010100111110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110110010100111111) && ({row_reg, col_reg}<19'b0110110010101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110010101000010) && ({row_reg, col_reg}<19'b0110110010101000101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110010101000101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110010101000110)) color_data = 12'b001001000010;
		if(({row_reg, col_reg}==19'b0110110010101000111)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0110110010101001000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110110010101001001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110010101001010) && ({row_reg, col_reg}<19'b0110110010101001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010101001100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110010101001101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0110110010101001110)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110110010101001111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110110010101010000) && ({row_reg, col_reg}<19'b0110110010101010010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110010101010010)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110010101010011)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==19'b0110110010101010100)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==19'b0110110010101010101)) color_data = 12'b001101010101;
		if(({row_reg, col_reg}==19'b0110110010101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010101010111)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110110010101011000)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110110010101011001)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0110110010101011010)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0110110010101011011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110110010101011100) && ({row_reg, col_reg}<19'b0110110010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110010101111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110110010101111001) && ({row_reg, col_reg}<19'b0110110010110110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110010110110100) && ({row_reg, col_reg}<19'b0110110010110111100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110110010110111100) && ({row_reg, col_reg}<19'b0110110011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110011001010001) && ({row_reg, col_reg}<19'b0110110011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110110011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110110011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110110100000000000) && ({row_reg, col_reg}<19'b0110110100010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100010100000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0110110100010100001) && ({row_reg, col_reg}<19'b0110110100010101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110110100010101001) && ({row_reg, col_reg}<19'b0110110100010101101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110110100010101101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0110110100010101110) && ({row_reg, col_reg}<19'b0110110100010110000)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0110110100010110000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110110100010110001)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0110110100010110010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=19'b0110110100010110011) && ({row_reg, col_reg}<19'b0110110100010110101)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==19'b0110110100010110101)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0110110100010110110)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0110110100010110111) && ({row_reg, col_reg}<19'b0110110100010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110110100010111111) && ({row_reg, col_reg}<19'b0110110100011010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100011010001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110110100011010010)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0110110100011010011) && ({row_reg, col_reg}<19'b0110110100011010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110100011010110)) color_data = 12'b010000110000;
		if(({row_reg, col_reg}>=19'b0110110100011010111) && ({row_reg, col_reg}<19'b0110110100011011001)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==19'b0110110100011011001)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==19'b0110110100011011010)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=19'b0110110100011011011) && ({row_reg, col_reg}<19'b0110110100011011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110100011011110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110110100011011111) && ({row_reg, col_reg}<19'b0110110100011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110100011110001) && ({row_reg, col_reg}<19'b0110110100011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110100011110011) && ({row_reg, col_reg}<19'b0110110100011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110110100011110110)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==19'b0110110100011110111)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==19'b0110110100011111000)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==19'b0110110100011111001)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0110110100011111010)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==19'b0110110100011111011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==19'b0110110100011111100)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110110100011111101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110100011111110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110100011111111)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}==19'b0110110100100000000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110100100000001) && ({row_reg, col_reg}<19'b0110110100100000011)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}>=19'b0110110100100000011) && ({row_reg, col_reg}<19'b0110110100100000101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110100100000101) && ({row_reg, col_reg}<19'b0110110100100000111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110100100000111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110100100001000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110100100001001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110100100001010)) color_data = 12'b001101010101;
		if(({row_reg, col_reg}==19'b0110110100100001011)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==19'b0110110100100001100)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==19'b0110110100100001101)) color_data = 12'b000100110011;
		if(({row_reg, col_reg}==19'b0110110100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100100001111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110100100010000) && ({row_reg, col_reg}<19'b0110110100100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100100011010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110100100011011)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110110100100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110110100100011101)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110110100100011110) && ({row_reg, col_reg}<19'b0110110100100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110100100100000) && ({row_reg, col_reg}<19'b0110110100100100110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110100100100110) && ({row_reg, col_reg}<19'b0110110100100101000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0110110100100101000) && ({row_reg, col_reg}<19'b0110110100100101011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110100100101011)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110110100100101100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110100100101101)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110110100100101110)) color_data = 12'b010001110100;
		if(({row_reg, col_reg}==19'b0110110100100101111)) color_data = 12'b101011001010;
		if(({row_reg, col_reg}==19'b0110110100100110000)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=19'b0110110100100110001) && ({row_reg, col_reg}<19'b0110110100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100100110011)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0110110100100110100) && ({row_reg, col_reg}<19'b0110110100100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100100110110)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0110110100100110111) && ({row_reg, col_reg}<19'b0110110100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100100111001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110110100100111010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110110100100111011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110110100100111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110100100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100100111110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110110100100111111) && ({row_reg, col_reg}<19'b0110110100101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100101000001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110100101000010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0110110100101000011) && ({row_reg, col_reg}<19'b0110110100101000101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110100101000101)) color_data = 12'b000100110001;
		if(({row_reg, col_reg}==19'b0110110100101000110)) color_data = 12'b011010000110;
		if(({row_reg, col_reg}==19'b0110110100101000111)) color_data = 12'b101011001010;
		if(({row_reg, col_reg}==19'b0110110100101001000)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0110110100101001001)) color_data = 12'b001001000010;
		if(({row_reg, col_reg}==19'b0110110100101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100101001011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110100101001100)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}>=19'b0110110100101001101) && ({row_reg, col_reg}<19'b0110110100101001111)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0110110100101001111)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==19'b0110110100101010000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110100101010001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110100101010010)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110100101010011)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==19'b0110110100101010100)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==19'b0110110100101010101)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0110110100101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100101010111)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110110100101011000)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0110110100101011001)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==19'b0110110100101011010)) color_data = 12'b010001100101;
		if(({row_reg, col_reg}==19'b0110110100101011011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110110100101011100) && ({row_reg, col_reg}<19'b0110110100101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100101011110)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}==19'b0110110100101011111)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==19'b0110110100101100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110110100101100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110100101100010) && ({row_reg, col_reg}<19'b0110110100101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110100101101000) && ({row_reg, col_reg}<19'b0110110100101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110100101111001) && ({row_reg, col_reg}<19'b0110110100101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110100101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110100101111110) && ({row_reg, col_reg}<19'b0110110100110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110100110110110) && ({row_reg, col_reg}<19'b0110110100110111010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110110100110111010) && ({row_reg, col_reg}<19'b0110110101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110101001010001) && ({row_reg, col_reg}<19'b0110110101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110110101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110110101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110110110000000000) && ({row_reg, col_reg}<19'b0110110110010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110110010100000) && ({row_reg, col_reg}<19'b0110110110010101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110110110010101000) && ({row_reg, col_reg}<19'b0110110110010101010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110110110010101010)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0110110110010101011) && ({row_reg, col_reg}<19'b0110110110010101101)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0110110110010101101) && ({row_reg, col_reg}<19'b0110110110010110000)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}>=19'b0110110110010110000) && ({row_reg, col_reg}<19'b0110110110010111000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110110110010111000) && ({row_reg, col_reg}<19'b0110110110010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110110110010111111) && ({row_reg, col_reg}<19'b0110110110011010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110110011010001) && ({row_reg, col_reg}<19'b0110110110011010011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110110110011010011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110110011010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110011010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110110011010110)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==19'b0110110110011010111)) color_data = 12'b010101000001;
		if(({row_reg, col_reg}==19'b0110110110011011000)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==19'b0110110110011011001)) color_data = 12'b010000110000;
		if(({row_reg, col_reg}==19'b0110110110011011010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=19'b0110110110011011011) && ({row_reg, col_reg}<19'b0110110110011011110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110110110011011110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110110110011011111) && ({row_reg, col_reg}<19'b0110110110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110110110011110001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==19'b0110110110011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110110011110011) && ({row_reg, col_reg}<19'b0110110110011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110011110110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110110011110111)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110110110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110011111001)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110110110011111010)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==19'b0110110110011111011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==19'b0110110110011111100)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==19'b0110110110011111101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110110011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110011111111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110100000001)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110110100000010)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}>=19'b0110110110100000011) && ({row_reg, col_reg}<19'b0110110110100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110100000101)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0110110110100000110)) color_data = 12'b000100110011;
		if(({row_reg, col_reg}==19'b0110110110100000111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110110110100001000) && ({row_reg, col_reg}<19'b0110110110100001010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110110100001010)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0110110110100001011)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==19'b0110110110100001100)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0110110110100001101)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110110110100001110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110110100001111)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}>=19'b0110110110100010000) && ({row_reg, col_reg}<19'b0110110110100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110100011001)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110110110100011010)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==19'b0110110110100011011)) color_data = 12'b010101100101;
		if(({row_reg, col_reg}==19'b0110110110100011100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==19'b0110110110100011101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==19'b0110110110100011110)) color_data = 12'b010101100101;
		if(({row_reg, col_reg}==19'b0110110110100011111)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110110110100100000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110110100100001)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110110110100100010)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0110110110100100011)) color_data = 12'b000100110000;
		if(({row_reg, col_reg}==19'b0110110110100100100)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0110110110100100101)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0110110110100100110)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0110110110100100111)) color_data = 12'b010101110100;
		if(({row_reg, col_reg}==19'b0110110110100101000)) color_data = 12'b001001000001;
		if(({row_reg, col_reg}>=19'b0110110110100101001) && ({row_reg, col_reg}<19'b0110110110100101011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110110100101011)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}>=19'b0110110110100101100) && ({row_reg, col_reg}<19'b0110110110100101110)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0110110110100101110)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0110110110100101111)) color_data = 12'b101111011010;
		if(({row_reg, col_reg}==19'b0110110110100110000)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==19'b0110110110100110001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110110100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110100110011)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0110110110100110100) && ({row_reg, col_reg}<19'b0110110110100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110100110110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110110110100110111) && ({row_reg, col_reg}<19'b0110110110100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110100111001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110110110100111010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110110110100111011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110110110100111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110110100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110100111110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110110110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110101000000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110110110101000001) && ({row_reg, col_reg}<19'b0110110110101000100)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110110110101000100)) color_data = 12'b000100110001;
		if(({row_reg, col_reg}==19'b0110110110101000101)) color_data = 12'b010001100100;
		if(({row_reg, col_reg}==19'b0110110110101000110)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0110110110101000111)) color_data = 12'b101011001010;
		if(({row_reg, col_reg}==19'b0110110110101001000)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0110110110101001001)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0110110110101001010)) color_data = 12'b000100110001;
		if(({row_reg, col_reg}==19'b0110110110101001011)) color_data = 12'b001101010011;
		if(({row_reg, col_reg}==19'b0110110110101001100)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0110110110101001101)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0110110110101001110)) color_data = 12'b101011011011;
		if(({row_reg, col_reg}==19'b0110110110101001111)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}>=19'b0110110110101010000) && ({row_reg, col_reg}<19'b0110110110101010011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110110110101010011)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==19'b0110110110101010100)) color_data = 12'b101011001100;
		if(({row_reg, col_reg}==19'b0110110110101010101)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0110110110101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110101010111)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110110110101011000)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0110110110101011001)) color_data = 12'b000101000011;
		if(({row_reg, col_reg}==19'b0110110110101011010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110110110101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110101011100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110110110101011101)) color_data = 12'b000101000011;
		if(({row_reg, col_reg}==19'b0110110110101011110)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0110110110101011111)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==19'b0110110110101100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110110110101100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0110110110101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110110101100011) && ({row_reg, col_reg}<19'b0110110110101100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110101100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110110101101000) && ({row_reg, col_reg}<19'b0110110110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110110110101111001) && ({row_reg, col_reg}<19'b0110110110101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110110110101111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110110110101111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110110110101111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0110110110101111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110110110110000000) && ({row_reg, col_reg}<19'b0110110111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110110111001010001) && ({row_reg, col_reg}<19'b0110110111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110110111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110110111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110111000000000000) && ({row_reg, col_reg}<19'b0110111000010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111000010100001) && ({row_reg, col_reg}<19'b0110111000010100100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110111000010100100)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0110111000010100101) && ({row_reg, col_reg}<19'b0110111000010101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110111000010101000) && ({row_reg, col_reg}<19'b0110111000010110000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110111000010110000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0110111000010110001)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0110111000010110010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110111000010110011) && ({row_reg, col_reg}<19'b0110111000010110101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110111000010110101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110111000010110110)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0110111000010110111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=19'b0110111000010111000) && ({row_reg, col_reg}<19'b0110111000010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110111000010111111) && ({row_reg, col_reg}<19'b0110111000011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111000011010000) && ({row_reg, col_reg}<19'b0110111000011010010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110111000011010010) && ({row_reg, col_reg}<19'b0110111000011010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110111000011010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000011010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110111000011010110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=19'b0110111000011010111) && ({row_reg, col_reg}<19'b0110111000011011001)) color_data = 12'b001100110000;
		if(({row_reg, col_reg}==19'b0110111000011011001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0110111000011011010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110111000011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111000011011100) && ({row_reg, col_reg}<19'b0110111000011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110111000011011111) && ({row_reg, col_reg}<19'b0110111000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111000011110000) && ({row_reg, col_reg}<19'b0110111000011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110111000011110011) && ({row_reg, col_reg}<19'b0110111000011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000011111010)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==19'b0110111000011111011)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0110111000011111100)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0110111000011111101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111000011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000011111111)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0110111000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000100000001)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0110111000100000010)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110111000100000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111000100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111000100000101) && ({row_reg, col_reg}<19'b0110111000100001000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111000100001000)) color_data = 12'b001101010101;
		if(({row_reg, col_reg}==19'b0110111000100001001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110111000100001010)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==19'b0110111000100001011)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0110111000100001100)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0110111000100001101)) color_data = 12'b000100110011;
		if(({row_reg, col_reg}==19'b0110111000100001110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111000100001111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110111000100010000) && ({row_reg, col_reg}<19'b0110111000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000100011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111000100011001)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==19'b0110111000100011010)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==19'b0110111000100011011)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==19'b0110111000100011100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110111000100011101)) color_data = 12'b101111001100;
		if(({row_reg, col_reg}==19'b0110111000100011110)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0110111000100011111)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==19'b0110111000100100000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110111000100100001)) color_data = 12'b000101000000;
		if(({row_reg, col_reg}==19'b0110111000100100010)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0110111000100100011)) color_data = 12'b010101110100;
		if(({row_reg, col_reg}==19'b0110111000100100100)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0110111000100100101)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0110111000100100110)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0110111000100100111)) color_data = 12'b101011001001;
		if(({row_reg, col_reg}==19'b0110111000100101000)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0110111000100101001)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0110111000100101010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111000100101011)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0110111000100101100)) color_data = 12'b100010110111;
		if(({row_reg, col_reg}>=19'b0110111000100101101) && ({row_reg, col_reg}<19'b0110111000100101111)) color_data = 12'b100010100111;
		if(({row_reg, col_reg}==19'b0110111000100101111)) color_data = 12'b101011001010;
		if(({row_reg, col_reg}==19'b0110111000100110000)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0110111000100110001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110111000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000100110011)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0110111000100110100) && ({row_reg, col_reg}<19'b0110111000100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000100110110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110111000100110111) && ({row_reg, col_reg}<19'b0110111000100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000100111001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110111000100111010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110111000100111011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110111000100111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110111000100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000100111110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110111000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000101000000)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}>=19'b0110111000101000001) && ({row_reg, col_reg}<19'b0110111000101000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111000101000011)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0110111000101000100)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}>=19'b0110111000101000101) && ({row_reg, col_reg}<19'b0110111000101000111)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0110111000101000111)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0110111000101001000)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0110111000101001001)) color_data = 12'b011010000110;
		if(({row_reg, col_reg}==19'b0110111000101001010)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0110111000101001011)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0110111000101001100)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0110111000101001101)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0110111000101001110)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0110111000101001111)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0110111000101010000)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}>=19'b0110111000101010001) && ({row_reg, col_reg}<19'b0110111000101010011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111000101010011)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0110111000101010100)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==19'b0110111000101010101)) color_data = 12'b001101010101;
		if(({row_reg, col_reg}==19'b0110111000101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000101010111)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0110111000101011000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111000101011001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111000101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000101011011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111000101011100)) color_data = 12'b000101000011;
		if(({row_reg, col_reg}==19'b0110111000101011101)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110111000101011110)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==19'b0110111000101011111)) color_data = 12'b110011101101;
		if(({row_reg, col_reg}==19'b0110111000101100000)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==19'b0110111000101100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111000101100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110111000101100011) && ({row_reg, col_reg}<19'b0110111000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000101111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110111000101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110111000101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111000101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110111000101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111000101111101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0110111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111000101111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0110111000110000000) && ({row_reg, col_reg}<19'b0110111001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111001001010001) && ({row_reg, col_reg}<19'b0110111001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110111001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110111001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110111010000000000) && ({row_reg, col_reg}<19'b0110111010010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111010010100001) && ({row_reg, col_reg}<19'b0110111010010100011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110111010010100011)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0110111010010100100) && ({row_reg, col_reg}<19'b0110111010010100110)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0110111010010100110) && ({row_reg, col_reg}<19'b0110111010010101000)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0110111010010101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110111010010101001) && ({row_reg, col_reg}<19'b0110111010010101100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110111010010101100) && ({row_reg, col_reg}<19'b0110111010010101110)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0110111010010101110) && ({row_reg, col_reg}<19'b0110111010010110000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0110111010010110000)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0110111010010110001)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0110111010010110010) && ({row_reg, col_reg}<19'b0110111010010110110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110111010010110110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0110111010010110111)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}>=19'b0110111010010111000) && ({row_reg, col_reg}<19'b0110111010010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110111010010111111) && ({row_reg, col_reg}<19'b0110111010011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111010011010000) && ({row_reg, col_reg}<19'b0110111010011010010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110111010011010010) && ({row_reg, col_reg}<19'b0110111010011010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110111010011010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111010011010101) && ({row_reg, col_reg}<19'b0110111010011010111)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0110111010011010111)) color_data = 12'b000100100000;
		if(({row_reg, col_reg}==19'b0110111010011011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0110111010011011001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0110111010011011010) && ({row_reg, col_reg}<19'b0110111010011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111010011011100) && ({row_reg, col_reg}<19'b0110111010011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110111010011011111) && ({row_reg, col_reg}<19'b0110111010011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111010011110010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110111010011110011) && ({row_reg, col_reg}<19'b0110111010011110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0110111010011110110) && ({row_reg, col_reg}<19'b0110111010011111000)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110111010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111010011111001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111010011111010)) color_data = 12'b010001100101;
		if(({row_reg, col_reg}==19'b0110111010011111011)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0110111010011111100)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==19'b0110111010011111101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111010011111111)) color_data = 12'b000101000011;
		if(({row_reg, col_reg}>=19'b0110111010100000000) && ({row_reg, col_reg}<19'b0110111010100000010)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0110111010100000010)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==19'b0110111010100000011)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110111010100000100)) color_data = 12'b001001010100;
		if(({row_reg, col_reg}>=19'b0110111010100000101) && ({row_reg, col_reg}<19'b0110111010100000111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111010100000111)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110111010100001000)) color_data = 12'b101011001100;
		if(({row_reg, col_reg}>=19'b0110111010100001001) && ({row_reg, col_reg}<19'b0110111010100001011)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0110111010100001011)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==19'b0110111010100001100)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0110111010100001101)) color_data = 12'b001001010100;
		if(({row_reg, col_reg}>=19'b0110111010100001110) && ({row_reg, col_reg}<19'b0110111010100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111010100011001)) color_data = 12'b010001100101;
		if(({row_reg, col_reg}==19'b0110111010100011010)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0110111010100011011)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==19'b0110111010100011100)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0110111010100011101)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0110111010100011110)) color_data = 12'b101111001100;
		if(({row_reg, col_reg}==19'b0110111010100011111)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==19'b0110111010100100000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110111010100100001)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0110111010100100010)) color_data = 12'b011010010101;
		if(({row_reg, col_reg}>=19'b0110111010100100011) && ({row_reg, col_reg}<19'b0110111010100100101)) color_data = 12'b100010110111;
		if(({row_reg, col_reg}==19'b0110111010100100101)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0110111010100100110)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0110111010100100111)) color_data = 12'b101111101010;
		if(({row_reg, col_reg}==19'b0110111010100101000)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0110111010100101001)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==19'b0110111010100101010)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0110111010100101011)) color_data = 12'b011010010101;
		if(({row_reg, col_reg}==19'b0110111010100101100)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0110111010100101101)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0110111010100101110)) color_data = 12'b011110100110;
		if(({row_reg, col_reg}==19'b0110111010100101111)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0110111010100110000)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==19'b0110111010100110001)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110111010100110010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111010100110011)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0110111010100110100) && ({row_reg, col_reg}<19'b0110111010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111010100110110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110111010100110111) && ({row_reg, col_reg}<19'b0110111010100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111010100111001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110111010100111010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110111010100111011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110111010100111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110111010100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111010100111110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110111010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111010101000000)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}>=19'b0110111010101000001) && ({row_reg, col_reg}<19'b0110111010101000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111010101000011)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0110111010101000100)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0110111010101000101)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0110111010101000110)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0110111010101000111)) color_data = 12'b001101100100;
		if(({row_reg, col_reg}==19'b0110111010101001000)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0110111010101001001)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0110111010101001010)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}>=19'b0110111010101001011) && ({row_reg, col_reg}<19'b0110111010101001101)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0110111010101001101)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0110111010101001110)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0110111010101001111)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}>=19'b0110111010101010000) && ({row_reg, col_reg}<19'b0110111010101010011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111010101010011)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110111010101010100)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==19'b0110111010101010101)) color_data = 12'b001101100101;
		if(({row_reg, col_reg}==19'b0110111010101010110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111010101010111)) color_data = 12'b010001100110;
		if(({row_reg, col_reg}==19'b0110111010101011000)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110111010101011001)) color_data = 12'b001001010100;
		if(({row_reg, col_reg}==19'b0110111010101011010)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111010101011011)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0110111010101011100)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==19'b0110111010101011101)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}>=19'b0110111010101011110) && ({row_reg, col_reg}<19'b0110111010101100000)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0110111010101100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111010101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111010101100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0110111010101100011) && ({row_reg, col_reg}<19'b0110111010101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111010101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0110111010101111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111010101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111010101111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111010101111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0110111010110000000) && ({row_reg, col_reg}<19'b0110111011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111011001010001) && ({row_reg, col_reg}<19'b0110111011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110111011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110111011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110111100000000000) && ({row_reg, col_reg}<19'b0110111100010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111100010100000) && ({row_reg, col_reg}<19'b0110111100010100101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110111100010100101) && ({row_reg, col_reg}<19'b0110111100010100111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110111100010100111)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0110111100010101000) && ({row_reg, col_reg}<19'b0110111100010101011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110111100010101011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0110111100010101100)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0110111100010101101) && ({row_reg, col_reg}<19'b0110111100010101111)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0110111100010101111)) color_data = 12'b001100000011;
		if(({row_reg, col_reg}==19'b0110111100010110000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0110111100010110001) && ({row_reg, col_reg}<19'b0110111100010110111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110111100010110111)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}>=19'b0110111100010111000) && ({row_reg, col_reg}<19'b0110111100010111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110111100010111111) && ({row_reg, col_reg}<19'b0110111100011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111100011010000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0110111100011010001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110111100011010010) && ({row_reg, col_reg}<19'b0110111100011010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110111100011010101) && ({row_reg, col_reg}<19'b0110111100011011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111100011011000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0110111100011011001) && ({row_reg, col_reg}<19'b0110111100011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111100011011100) && ({row_reg, col_reg}<19'b0110111100011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110111100011011111) && ({row_reg, col_reg}<19'b0110111100011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111100011110011) && ({row_reg, col_reg}<19'b0110111100011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110111100011110101)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0110111100011110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110111100011110111)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110111100011111000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110111100011111001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111100011111010)) color_data = 12'b001001000100;
		if(({row_reg, col_reg}==19'b0110111100011111011)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0110111100011111100)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0110111100011111101)) color_data = 12'b000100110011;
		if(({row_reg, col_reg}==19'b0110111100011111110)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111100011111111)) color_data = 12'b001101100101;
		if(({row_reg, col_reg}==19'b0110111100100000000)) color_data = 12'b110011111110;
		if(({row_reg, col_reg}>=19'b0110111100100000001) && ({row_reg, col_reg}<19'b0110111100100000011)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0110111100100000011)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==19'b0110111100100000100)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}>=19'b0110111100100000101) && ({row_reg, col_reg}<19'b0110111100100000111)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0110111100100000111)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0110111100100001000)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==19'b0110111100100001001)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0110111100100001010)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==19'b0110111100100001011)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0110111100100001100)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0110111100100001101)) color_data = 12'b001101100101;
		if(({row_reg, col_reg}==19'b0110111100100001110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110111100100001111) && ({row_reg, col_reg}<19'b0110111100100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111100100011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111100100011001)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0110111100100011010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110111100100011011)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==19'b0110111100100011100)) color_data = 12'b010001100101;
		if(({row_reg, col_reg}==19'b0110111100100011101)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110111100100011110)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0110111100100011111)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0110111100100100000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111100100100001)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0110111100100100010)) color_data = 12'b011110100110;
		if(({row_reg, col_reg}==19'b0110111100100100011)) color_data = 12'b100011001000;
		if(({row_reg, col_reg}==19'b0110111100100100100)) color_data = 12'b100010110111;
		if(({row_reg, col_reg}>=19'b0110111100100100101) && ({row_reg, col_reg}<19'b0110111100100100111)) color_data = 12'b011010100110;
		if(({row_reg, col_reg}==19'b0110111100100100111)) color_data = 12'b011110100110;
		if(({row_reg, col_reg}==19'b0110111100100101000)) color_data = 12'b100111011001;
		if(({row_reg, col_reg}==19'b0110111100100101001)) color_data = 12'b001101110011;
		if(({row_reg, col_reg}==19'b0110111100100101010)) color_data = 12'b001001100010;
		if(({row_reg, col_reg}==19'b0110111100100101011)) color_data = 12'b100010110111;
		if(({row_reg, col_reg}==19'b0110111100100101100)) color_data = 12'b100111001000;
		if(({row_reg, col_reg}>=19'b0110111100100101101) && ({row_reg, col_reg}<19'b0110111100100101111)) color_data = 12'b010001110011;
		if(({row_reg, col_reg}==19'b0110111100100101111)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0110111100100110000)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==19'b0110111100100110001)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110111100100110010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111100100110011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110111100100110100) && ({row_reg, col_reg}<19'b0110111100100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111100100110110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}>=19'b0110111100100110111) && ({row_reg, col_reg}<19'b0110111100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111100100111001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110111100100111010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110111100100111011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110111100100111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110111100100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111100100111110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110111100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111100101000000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110111100101000001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111100101000010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110111100101000011)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0110111100101000100)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0110111100101000101)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0110111100101000110)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0110111100101000111)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0110111100101001000)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0110111100101001001)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0110111100101001010)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0110111100101001011)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0110111100101001100)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0110111100101001101)) color_data = 12'b010001110100;
		if(({row_reg, col_reg}==19'b0110111100101001110)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0110111100101001111)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0110111100101010000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111100101010001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111100101010010)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111100101010011)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110111100101010100)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==19'b0110111100101010101)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==19'b0110111100101010110)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111100101010111)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110111100101011000)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==19'b0110111100101011001)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}>=19'b0110111100101011010) && ({row_reg, col_reg}<19'b0110111100101011100)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0110111100101011100)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}>=19'b0110111100101011101) && ({row_reg, col_reg}<19'b0110111100101011111)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==19'b0110111100101011111)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0110111100101100000)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==19'b0110111100101100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0110111100101100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110111100101100011) && ({row_reg, col_reg}<19'b0110111100101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111100101111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110111100101111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111100101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111100101111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0110111100110000000) && ({row_reg, col_reg}<19'b0110111101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111101001010001) && ({row_reg, col_reg}<19'b0110111101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110111101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110111101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0110111110000000000) && ({row_reg, col_reg}<19'b0110111110010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110010100000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110111110010100001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0110111110010100010) && ({row_reg, col_reg}<19'b0110111110010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111110010100111) && ({row_reg, col_reg}<19'b0110111110010101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110111110010101001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0110111110010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111110010101011) && ({row_reg, col_reg}<19'b0110111110010110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110111110010110000) && ({row_reg, col_reg}<19'b0110111110010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111110010110010) && ({row_reg, col_reg}<19'b0110111110010110110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0110111110010110110) && ({row_reg, col_reg}<19'b0110111110011010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110011010000)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0110111110011010001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0110111110011010010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110111110011010011) && ({row_reg, col_reg}<19'b0110111110011010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110011010101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110111110011010110) && ({row_reg, col_reg}<19'b0110111110011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110011011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110111110011011001) && ({row_reg, col_reg}<19'b0110111110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111110011011101) && ({row_reg, col_reg}<19'b0110111110011011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0110111110011011111) && ({row_reg, col_reg}<19'b0110111110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110011111000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110111110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110011111010)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111110011111011)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==19'b0110111110011111100)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0110111110011111101)) color_data = 12'b001001010100;
		if(({row_reg, col_reg}==19'b0110111110011111110)) color_data = 12'b000101000011;
		if(({row_reg, col_reg}==19'b0110111110011111111)) color_data = 12'b010110010111;
		if(({row_reg, col_reg}==19'b0110111110100000000)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==19'b0110111110100000001)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0110111110100000010)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0110111110100000011)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==19'b0110111110100000100)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==19'b0110111110100000101)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110111110100000110)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0110111110100000111)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0110111110100001000)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0110111110100001001)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0110111110100001010)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0110111110100001011)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0110111110100001100)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0110111110100001101)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0110111110100001110)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0110111110100001111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0110111110100010000) && ({row_reg, col_reg}<19'b0110111110100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110100011000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110111110100011001)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==19'b0110111110100011010)) color_data = 12'b101011001100;
		if(({row_reg, col_reg}==19'b0110111110100011011)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==19'b0110111110100011100)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110111110100011101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==19'b0110111110100011110)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==19'b0110111110100011111)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0110111110100100000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111110100100001)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==19'b0110111110100100010)) color_data = 12'b011010100110;
		if(({row_reg, col_reg}==19'b0110111110100100011)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0110111110100100100)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0110111110100100101)) color_data = 12'b010001110011;
		if(({row_reg, col_reg}==19'b0110111110100100110)) color_data = 12'b001101100010;
		if(({row_reg, col_reg}==19'b0110111110100100111)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0110111110100101000)) color_data = 12'b011110110111;
		if(({row_reg, col_reg}==19'b0110111110100101001)) color_data = 12'b001101110011;
		if(({row_reg, col_reg}==19'b0110111110100101010)) color_data = 12'b010010000100;
		if(({row_reg, col_reg}==19'b0110111110100101011)) color_data = 12'b100011001000;
		if(({row_reg, col_reg}==19'b0110111110100101100)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0110111110100101101)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0110111110100101110)) color_data = 12'b000001000000;
		if(({row_reg, col_reg}==19'b0110111110100101111)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0110111110100110000)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0110111110100110001)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0110111110100110010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111110100110011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0110111110100110100) && ({row_reg, col_reg}<19'b0110111110100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110100110110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110111110100110111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111110100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110100111001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0110111110100111010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==19'b0110111110100111011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0110111110100111100)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0110111110100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110100111110)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0110111110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110101000000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111110101000001)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110111110101000010)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0110111110101000011)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0110111110101000100)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0110111110101000101)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0110111110101000110)) color_data = 12'b100111011010;
		if(({row_reg, col_reg}==19'b0110111110101000111)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0110111110101001000)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0110111110101001001)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110111110101001010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111110101001011)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0110111110101001100)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0110111110101001101)) color_data = 12'b100011001001;
		if(({row_reg, col_reg}==19'b0110111110101001110)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0110111110101001111)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0110111110101010000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0110111110101010001) && ({row_reg, col_reg}<19'b0110111110101010011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111110101010011)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0110111110101010100)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==19'b0110111110101010101)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==19'b0110111110101010110)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0110111110101010111)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0110111110101011000)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==19'b0110111110101011001)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0110111110101011010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0110111110101011011)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0110111110101011100)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0110111110101011101)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==19'b0110111110101011110)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==19'b0110111110101011111)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==19'b0110111110101100000)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==19'b0110111110101100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0110111110101100010) && ({row_reg, col_reg}<19'b0110111110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0110111110101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0110111110101111001)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0110111110101111010)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==19'b0110111110101111011)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==19'b0110111110101111100)) color_data = 12'b110111011011;
		if(({row_reg, col_reg}==19'b0110111110101111101)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==19'b0110111110101111110)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==19'b0110111110101111111)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}>=19'b0110111110110000000) && ({row_reg, col_reg}<19'b0110111111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0110111111001010001) && ({row_reg, col_reg}<19'b0110111111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0110111111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0110111111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111000000000000000) && ({row_reg, col_reg}<19'b0111000000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000011110000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111000000011110001) && ({row_reg, col_reg}<19'b0111000000011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000011110011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000000011110100)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000000011110101)) color_data = 12'b000000100010;
		if(({row_reg, col_reg}==19'b0111000000011110110)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000000011110111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000000011111000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000000011111001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000000011111010)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0111000000011111011)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0111000000011111100)) color_data = 12'b100011001011;
		if(({row_reg, col_reg}==19'b0111000000011111101)) color_data = 12'b001101110101;
		if(({row_reg, col_reg}==19'b0111000000011111110)) color_data = 12'b001101110110;
		if(({row_reg, col_reg}==19'b0111000000011111111)) color_data = 12'b100111011100;
		if(({row_reg, col_reg}==19'b0111000000100000000)) color_data = 12'b001001100011;
		if(({row_reg, col_reg}==19'b0111000000100000001)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0111000000100000010)) color_data = 12'b010001110100;
		if(({row_reg, col_reg}==19'b0111000000100000011)) color_data = 12'b100011001000;
		if(({row_reg, col_reg}==19'b0111000000100000100)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0111000000100000101)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0111000000100000110)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0111000000100000111)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111000000100001000)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0111000000100001001)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111000000100001010)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000000100001011)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0111000000100001100)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0111000000100001101)) color_data = 12'b010001110100;
		if(({row_reg, col_reg}>=19'b0111000000100001110) && ({row_reg, col_reg}<19'b0111000000100010000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0111000000100010000) && ({row_reg, col_reg}<19'b0111000000100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000100011000)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==19'b0111000000100011001)) color_data = 12'b010001100101;
		if(({row_reg, col_reg}==19'b0111000000100011010)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0111000000100011011)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0111000000100011100)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==19'b0111000000100011101)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0111000000100011110)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==19'b0111000000100011111)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0111000000100100000)) color_data = 12'b000100110001;
		if(({row_reg, col_reg}==19'b0111000000100100001)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000000100100010)) color_data = 12'b010001110100;
		if(({row_reg, col_reg}==19'b0111000000100100011)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0111000000100100100)) color_data = 12'b011110111000;
		if(({row_reg, col_reg}>=19'b0111000000100100101) && ({row_reg, col_reg}<19'b0111000000100100111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000000100100111)) color_data = 12'b010110010110;
		if(({row_reg, col_reg}==19'b0111000000100101000)) color_data = 12'b011110111000;
		if(({row_reg, col_reg}>=19'b0111000000100101001) && ({row_reg, col_reg}<19'b0111000000100101011)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0111000000100101011)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111000000100101100)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0111000000100101101)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000000100101110)) color_data = 12'b010001110100;
		if(({row_reg, col_reg}==19'b0111000000100101111)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0111000000100110000)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000000100110001)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0111000000100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000100110011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000000100110100)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111000000100110101) && ({row_reg, col_reg}<19'b0111000000100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000100110111)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0111000000100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000100111001)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==19'b0111000000100111010)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==19'b0111000000100111011)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0111000000100111100)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}>=19'b0111000000100111101) && ({row_reg, col_reg}<19'b0111000000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000100111111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000000101000000)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000000101000001)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000000101000010)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000000101000011)) color_data = 12'b010001110100;
		if(({row_reg, col_reg}==19'b0111000000101000100)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000000101000101)) color_data = 12'b100111011010;
		if(({row_reg, col_reg}==19'b0111000000101000110)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0111000000101000111)) color_data = 12'b001101100100;
		if(({row_reg, col_reg}==19'b0111000000101001000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000000101001001)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0111000000101001010)) color_data = 12'b000001000001;
		if(({row_reg, col_reg}==19'b0111000000101001011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000000101001100)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000000101001101)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0111000000101001110)) color_data = 12'b110111111101;
		if(({row_reg, col_reg}==19'b0111000000101001111)) color_data = 12'b111011111110;
		if(({row_reg, col_reg}==19'b0111000000101010000)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111000000101010001)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000000101010010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000000101010011)) color_data = 12'b010110010110;
		if(({row_reg, col_reg}==19'b0111000000101010100)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0111000000101010101)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111000000101010110)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}==19'b0111000000101010111)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111000000101011000)) color_data = 12'b100111011010;
		if(({row_reg, col_reg}==19'b0111000000101011001)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0111000000101011010)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000000101011011)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0111000000101011100)) color_data = 12'b101011011011;
		if(({row_reg, col_reg}==19'b0111000000101011101)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111000000101011110)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0111000000101011111)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111000000101100000)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0111000000101100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111000000101100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111000000101100011) && ({row_reg, col_reg}<19'b0111000000101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000101100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111000000101100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111000000101100111) && ({row_reg, col_reg}<19'b0111000000101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000101110001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111000000101110010) && ({row_reg, col_reg}<19'b0111000000101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000101111001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0111000000101111010)) color_data = 12'b011110000100;
		if(({row_reg, col_reg}==19'b0111000000101111011)) color_data = 12'b101111001000;
		if(({row_reg, col_reg}>=19'b0111000000101111100) && ({row_reg, col_reg}<19'b0111000000101111110)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0111000000101111110)) color_data = 12'b110011011000;
		if(({row_reg, col_reg}==19'b0111000000101111111)) color_data = 12'b100010010100;
		if(({row_reg, col_reg}==19'b0111000000110000000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==19'b0111000000110000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111000000110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111000000110000011) && ({row_reg, col_reg}<19'b0111000000110000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000000110000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111000000110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111000000110000111) && ({row_reg, col_reg}<19'b0111000001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111000001001010001) && ({row_reg, col_reg}<19'b0111000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111000001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111000001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111000010000000000) && ({row_reg, col_reg}<19'b0111000010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000010011110000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111000010011110001) && ({row_reg, col_reg}<19'b0111000010011110011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111000010011110011) && ({row_reg, col_reg}<19'b0111000010011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000010011110101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000010011110110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111000010011110111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000010011111000)) color_data = 12'b001001010100;
		if(({row_reg, col_reg}==19'b0111000010011111001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000010011111010)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000010011111011)) color_data = 12'b011010101001;
		if(({row_reg, col_reg}==19'b0111000010011111100)) color_data = 12'b100011001011;
		if(({row_reg, col_reg}==19'b0111000010011111101)) color_data = 12'b010010000111;
		if(({row_reg, col_reg}==19'b0111000010011111110)) color_data = 12'b001110000110;
		if(({row_reg, col_reg}==19'b0111000010011111111)) color_data = 12'b100011001010;
		if(({row_reg, col_reg}==19'b0111000010100000000)) color_data = 12'b001101110011;
		if(({row_reg, col_reg}==19'b0111000010100000001)) color_data = 12'b001101100010;
		if(({row_reg, col_reg}==19'b0111000010100000010)) color_data = 12'b011010010101;
		if(({row_reg, col_reg}==19'b0111000010100000011)) color_data = 12'b101011011001;
		if(({row_reg, col_reg}==19'b0111000010100000100)) color_data = 12'b100011001000;
		if(({row_reg, col_reg}==19'b0111000010100000101)) color_data = 12'b001101110011;
		if(({row_reg, col_reg}==19'b0111000010100000110)) color_data = 12'b010001110011;
		if(({row_reg, col_reg}==19'b0111000010100000111)) color_data = 12'b100011001000;
		if(({row_reg, col_reg}==19'b0111000010100001000)) color_data = 12'b010001110011;
		if(({row_reg, col_reg}>=19'b0111000010100001001) && ({row_reg, col_reg}<19'b0111000010100001011)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000010100001011)) color_data = 12'b010110000100;
		if(({row_reg, col_reg}==19'b0111000010100001100)) color_data = 12'b100010110111;
		if(({row_reg, col_reg}==19'b0111000010100001101)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0111000010100001110)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000010100001111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111000010100010000) && ({row_reg, col_reg}<19'b0111000010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000010100011000)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0111000010100011001)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0111000010100011010)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==19'b0111000010100011011)) color_data = 12'b101111001100;
		if(({row_reg, col_reg}==19'b0111000010100011100)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==19'b0111000010100011101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==19'b0111000010100011110)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0111000010100011111)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0111000010100100000)) color_data = 12'b001001000010;
		if(({row_reg, col_reg}==19'b0111000010100100001)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0111000010100100010)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111000010100100011)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0111000010100100100)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}>=19'b0111000010100100101) && ({row_reg, col_reg}<19'b0111000010100100111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000010100100111)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111000010100101000)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000010100101001)) color_data = 12'b011110111000;
		if(({row_reg, col_reg}>=19'b0111000010100101010) && ({row_reg, col_reg}<19'b0111000010100101100)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111000010100101100)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0111000010100101101)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111000010100101110)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111000010100101111)) color_data = 12'b110011111100;
		if(({row_reg, col_reg}==19'b0111000010100110000)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111000010100110001)) color_data = 12'b000101000011;
		if(({row_reg, col_reg}==19'b0111000010100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000010100110011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000010100110100)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000010100110101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000010100110111)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0111000010100111000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000010100111001)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0111000010100111010)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==19'b0111000010100111011)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0111000010100111100)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}>=19'b0111000010100111101) && ({row_reg, col_reg}<19'b0111000010100111111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000010100111111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111000010101000000) && ({row_reg, col_reg}<19'b0111000010101000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000010101000011)) color_data = 12'b001001100011;
		if(({row_reg, col_reg}>=19'b0111000010101000100) && ({row_reg, col_reg}<19'b0111000010101000110)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0111000010101000110)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0111000010101000111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000010101001000)) color_data = 12'b001101100100;
		if(({row_reg, col_reg}>=19'b0111000010101001001) && ({row_reg, col_reg}<19'b0111000010101001011)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111000010101001011)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111000010101001100)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000010101001101)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}==19'b0111000010101001110)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111000010101001111)) color_data = 12'b011110111000;
		if(({row_reg, col_reg}==19'b0111000010101010000)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0111000010101010001)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111000010101010010)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000010101010011)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111000010101010100)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0111000010101010101)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111000010101010110)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111000010101010111)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000010101011000)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111000010101011001)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0111000010101011010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000010101011011)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000010101011100)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000010101011101)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0111000010101011110)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0111000010101011111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000010101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111000010101100001) && ({row_reg, col_reg}<19'b0111000010101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111000010101100011) && ({row_reg, col_reg}<19'b0111000010101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111000010101110000) && ({row_reg, col_reg}<19'b0111000010101110011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111000010101110011) && ({row_reg, col_reg}<19'b0111000010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000010101111000)) color_data = 12'b011001100011;
		if(({row_reg, col_reg}==19'b0111000010101111001)) color_data = 12'b101010110111;
		if(({row_reg, col_reg}==19'b0111000010101111010)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}>=19'b0111000010101111011) && ({row_reg, col_reg}<19'b0111000010101111101)) color_data = 12'b110111101000;
		if(({row_reg, col_reg}==19'b0111000010101111101)) color_data = 12'b110111111000;
		if(({row_reg, col_reg}==19'b0111000010101111110)) color_data = 12'b110111100111;
		if(({row_reg, col_reg}==19'b0111000010101111111)) color_data = 12'b110011011000;
		if(({row_reg, col_reg}==19'b0111000010110000000)) color_data = 12'b100110101000;
		if(({row_reg, col_reg}==19'b0111000010110000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111000010110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000010110000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111000010110000100) && ({row_reg, col_reg}<19'b0111000011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111000011001010001) && ({row_reg, col_reg}<19'b0111000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111000011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111000011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111000100000000000) && ({row_reg, col_reg}<19'b0111000100011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111000100011110001) && ({row_reg, col_reg}<19'b0111000100011110011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111000100011110011) && ({row_reg, col_reg}<19'b0111000100011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000100011110110)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000100011110111)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0111000100011111000)) color_data = 12'b001101100101;
		if(({row_reg, col_reg}>=19'b0111000100011111001) && ({row_reg, col_reg}<19'b0111000100011111011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000100011111011)) color_data = 12'b010010000110;
		if(({row_reg, col_reg}==19'b0111000100011111100)) color_data = 12'b011110111010;
		if(({row_reg, col_reg}==19'b0111000100011111101)) color_data = 12'b010110010111;
		if(({row_reg, col_reg}==19'b0111000100011111110)) color_data = 12'b010010000111;
		if(({row_reg, col_reg}==19'b0111000100011111111)) color_data = 12'b011110111001;
		if(({row_reg, col_reg}==19'b0111000100100000000)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111000100100000001)) color_data = 12'b010110000100;
		if(({row_reg, col_reg}==19'b0111000100100000010)) color_data = 12'b011110100111;
		if(({row_reg, col_reg}==19'b0111000100100000011)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0111000100100000100)) color_data = 12'b100111001000;
		if(({row_reg, col_reg}>=19'b0111000100100000101) && ({row_reg, col_reg}<19'b0111000100100000111)) color_data = 12'b010110000100;
		if(({row_reg, col_reg}==19'b0111000100100000111)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111000100100001000)) color_data = 12'b011010010101;
		if(({row_reg, col_reg}==19'b0111000100100001001)) color_data = 12'b001001010001;
		if(({row_reg, col_reg}==19'b0111000100100001010)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0111000100100001011)) color_data = 12'b011110100110;
		if(({row_reg, col_reg}==19'b0111000100100001100)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111000100100001101)) color_data = 12'b010001110011;
		if(({row_reg, col_reg}==19'b0111000100100001110)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000100100001111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111000100100010000) && ({row_reg, col_reg}<19'b0111000100100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000100100011000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0111000100100011001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0111000100100011010)) color_data = 12'b110111111110;
		if(({row_reg, col_reg}==19'b0111000100100011011)) color_data = 12'b110011011101;
		if(({row_reg, col_reg}==19'b0111000100100011100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==19'b0111000100100011101)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==19'b0111000100100011110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==19'b0111000100100011111)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0111000100100100000)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0111000100100100001)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}==19'b0111000100100100010)) color_data = 12'b010101110101;
		if(({row_reg, col_reg}==19'b0111000100100100011)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0111000100100100100)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}>=19'b0111000100100100101) && ({row_reg, col_reg}<19'b0111000100100100111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000100100100111)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0111000100100101000)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0111000100100101001)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111000100100101010)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0111000100100101011)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0111000100100101100)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111000100100101101)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000100100101110)) color_data = 12'b100110111001;
		if(({row_reg, col_reg}==19'b0111000100100101111)) color_data = 12'b101011011011;
		if(({row_reg, col_reg}==19'b0111000100100110000)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0111000100100110001)) color_data = 12'b001001010100;
		if(({row_reg, col_reg}==19'b0111000100100110010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111000100100110011) && ({row_reg, col_reg}<19'b0111000100100110101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111000100100110101) && ({row_reg, col_reg}<19'b0111000100100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000100100110111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000100100111000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000100100111001)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==19'b0111000100100111010)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0111000100100111011)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0111000100100111100)) color_data = 12'b000101000011;
		if(({row_reg, col_reg}==19'b0111000100100111101)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0111000100100111110)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0111000100100111111)) color_data = 12'b001101100100;
		if(({row_reg, col_reg}==19'b0111000100101000000)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}>=19'b0111000100101000001) && ({row_reg, col_reg}<19'b0111000100101000011)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111000100101000011)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0111000100101000100)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0111000100101000101)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0111000100101000110)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111000100101000111)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0111000100101001000)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111000100101001001)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000100101001010)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0111000100101001011)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0111000100101001100)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0111000100101001101)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000100101001110)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}==19'b0111000100101001111)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111000100101010000)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000100101010001)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0111000100101010010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000100101010011)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111000100101010100)) color_data = 12'b100111001001;
		if(({row_reg, col_reg}==19'b0111000100101010101)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0111000100101010110)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}==19'b0111000100101010111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000100101011000)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111000100101011001)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000100101011010)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0111000100101011011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000100101011100)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0111000100101011101)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0111000100101011110)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}>=19'b0111000100101011111) && ({row_reg, col_reg}<19'b0111000100101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000100101100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111000100101100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111000100101100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111000100101100100) && ({row_reg, col_reg}<19'b0111000100101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111000100101110000) && ({row_reg, col_reg}<19'b0111000100101110011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111000100101110011) && ({row_reg, col_reg}<19'b0111000100101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000100101111000)) color_data = 12'b100010000101;
		if(({row_reg, col_reg}==19'b0111000100101111001)) color_data = 12'b110111101010;
		if(({row_reg, col_reg}==19'b0111000100101111010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==19'b0111000100101111011)) color_data = 12'b111111111011;
		if(({row_reg, col_reg}==19'b0111000100101111100)) color_data = 12'b110111101000;
		if(({row_reg, col_reg}==19'b0111000100101111101)) color_data = 12'b110111100111;
		if(({row_reg, col_reg}==19'b0111000100101111110)) color_data = 12'b111011111000;
		if(({row_reg, col_reg}==19'b0111000100101111111)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==19'b0111000100110000000)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==19'b0111000100110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000100110000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111000100110000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111000100110000100) && ({row_reg, col_reg}<19'b0111000100110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000100110000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111000100110001000) && ({row_reg, col_reg}<19'b0111000101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111000101001010001) && ({row_reg, col_reg}<19'b0111000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111000101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111000101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111000110000000000) && ({row_reg, col_reg}<19'b0111000110011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000110011110001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000110011110010)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0111000110011110011) && ({row_reg, col_reg}<19'b0111000110011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000110011110110)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0111000110011110111)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==19'b0111000110011111000)) color_data = 12'b001101100101;
		if(({row_reg, col_reg}==19'b0111000110011111001)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000110011111010)) color_data = 12'b000000110010;
		if(({row_reg, col_reg}==19'b0111000110011111011)) color_data = 12'b010010000110;
		if(({row_reg, col_reg}==19'b0111000110011111100)) color_data = 12'b011010101000;
		if(({row_reg, col_reg}==19'b0111000110011111101)) color_data = 12'b010010000110;
		if(({row_reg, col_reg}==19'b0111000110011111110)) color_data = 12'b010010000111;
		if(({row_reg, col_reg}==19'b0111000110011111111)) color_data = 12'b100011001010;
		if(({row_reg, col_reg}==19'b0111000110100000000)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}>=19'b0111000110100000001) && ({row_reg, col_reg}<19'b0111000110100000011)) color_data = 12'b011110100110;
		if(({row_reg, col_reg}==19'b0111000110100000011)) color_data = 12'b100010110111;
		if(({row_reg, col_reg}==19'b0111000110100000100)) color_data = 12'b011010010110;
		if(({row_reg, col_reg}==19'b0111000110100000101)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0111000110100000110)) color_data = 12'b010001110011;
		if(({row_reg, col_reg}==19'b0111000110100000111)) color_data = 12'b011110100110;
		if(({row_reg, col_reg}==19'b0111000110100001000)) color_data = 12'b101111101011;
		if(({row_reg, col_reg}==19'b0111000110100001001)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111000110100001010)) color_data = 12'b100010110111;
		if(({row_reg, col_reg}>=19'b0111000110100001011) && ({row_reg, col_reg}<19'b0111000110100001101)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0111000110100001101)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111000110100001110)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111000110100001111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111000110100010000) && ({row_reg, col_reg}<19'b0111000110100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000110100011001)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==19'b0111000110100011010)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==19'b0111000110100011011)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0111000110100011100)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==19'b0111000110100011101)) color_data = 12'b001000110011;
		if(({row_reg, col_reg}==19'b0111000110100011110)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==19'b0111000110100011111)) color_data = 12'b110011101101;
		if(({row_reg, col_reg}==19'b0111000110100100000)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0111000110100100001)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}==19'b0111000110100100010)) color_data = 12'b001101100100;
		if(({row_reg, col_reg}==19'b0111000110100100011)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0111000110100100100)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}>=19'b0111000110100100101) && ({row_reg, col_reg}<19'b0111000110100100111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111000110100100111) && ({row_reg, col_reg}<19'b0111000110100101001)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0111000110100101001)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111000110100101010)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0111000110100101011)) color_data = 12'b011010000110;
		if(({row_reg, col_reg}==19'b0111000110100101100)) color_data = 12'b100010101000;
		if(({row_reg, col_reg}==19'b0111000110100101101)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0111000110100101110)) color_data = 12'b010101110101;
		if(({row_reg, col_reg}==19'b0111000110100101111)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0111000110100110000)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0111000110100110001)) color_data = 12'b000101000011;
		if(({row_reg, col_reg}==19'b0111000110100110010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111000110100110011) && ({row_reg, col_reg}<19'b0111000110100110101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111000110100110101) && ({row_reg, col_reg}<19'b0111000110100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000110100110111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111000110100111000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000110100111001)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==19'b0111000110100111010)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==19'b0111000110100111011)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0111000110100111100)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0111000110100111101)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==19'b0111000110100111110)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==19'b0111000110100111111)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0111000110101000000)) color_data = 12'b110011101100;
		if(({row_reg, col_reg}==19'b0111000110101000001)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0111000110101000010)) color_data = 12'b001101010011;
		if(({row_reg, col_reg}==19'b0111000110101000011)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}==19'b0111000110101000100)) color_data = 12'b001101100100;
		if(({row_reg, col_reg}==19'b0111000110101000101)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0111000110101000110)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111000110101000111)) color_data = 12'b101011011011;
		if(({row_reg, col_reg}==19'b0111000110101001000)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}>=19'b0111000110101001001) && ({row_reg, col_reg}<19'b0111000110101001011)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}>=19'b0111000110101001011) && ({row_reg, col_reg}<19'b0111000110101001101)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}>=19'b0111000110101001101) && ({row_reg, col_reg}<19'b0111000110101001111)) color_data = 12'b010101110101;
		if(({row_reg, col_reg}==19'b0111000110101001111)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111000110101010000)) color_data = 12'b100010101000;
		if(({row_reg, col_reg}==19'b0111000110101010001)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}==19'b0111000110101010010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111000110101010011)) color_data = 12'b001101100100;
		if(({row_reg, col_reg}==19'b0111000110101010100)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000110101010101)) color_data = 12'b011110101000;
		if(({row_reg, col_reg}==19'b0111000110101010110)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0111000110101010111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000110101011000)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==19'b0111000110101011001)) color_data = 12'b101111011011;
		if(({row_reg, col_reg}==19'b0111000110101011010)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0111000110101011011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111000110101011100)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111000110101011101)) color_data = 12'b101111101011;
		if(({row_reg, col_reg}==19'b0111000110101011110)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0111000110101011111)) color_data = 12'b000100110001;
		if(({row_reg, col_reg}==19'b0111000110101100000)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==19'b0111000110101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000110101100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111000110101100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111000110101100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111000110101100101) && ({row_reg, col_reg}<19'b0111000110101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111000110101110000) && ({row_reg, col_reg}<19'b0111000110101110010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111000110101110010) && ({row_reg, col_reg}<19'b0111000110101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000110101111001)) color_data = 12'b011001110011;
		if(({row_reg, col_reg}==19'b0111000110101111010)) color_data = 12'b110011011000;
		if(({row_reg, col_reg}>=19'b0111000110101111011) && ({row_reg, col_reg}<19'b0111000110101111101)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0111000110101111101)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}==19'b0111000110101111110)) color_data = 12'b110111101000;
		if(({row_reg, col_reg}==19'b0111000110101111111)) color_data = 12'b110011011000;
		if(({row_reg, col_reg}==19'b0111000110110000000)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==19'b0111000110110000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111000110110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000110110000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111000110110000100) && ({row_reg, col_reg}<19'b0111000110110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111000110110000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111000110110001000) && ({row_reg, col_reg}<19'b0111000111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111000111001010001) && ({row_reg, col_reg}<19'b0111000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111000111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111000111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111001000000000000) && ({row_reg, col_reg}<19'b0111001000011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000011110010)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0111001000011110011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001000011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000011110101)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001000011110110)) color_data = 12'b001101010101;
		if(({row_reg, col_reg}>=19'b0111001000011110111) && ({row_reg, col_reg}<19'b0111001000011111001)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0111001000011111001)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0111001000011111010)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0111001000011111011)) color_data = 12'b011110111001;
		if(({row_reg, col_reg}==19'b0111001000011111100)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0111001000011111101)) color_data = 12'b000101010011;
		if(({row_reg, col_reg}==19'b0111001000011111110)) color_data = 12'b001101110101;
		if(({row_reg, col_reg}==19'b0111001000011111111)) color_data = 12'b100011001010;
		if(({row_reg, col_reg}==19'b0111001000100000000)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0111001000100000001)) color_data = 12'b100010100111;
		if(({row_reg, col_reg}==19'b0111001000100000010)) color_data = 12'b010110000101;
		if(({row_reg, col_reg}==19'b0111001000100000011)) color_data = 12'b001101100011;
		if(({row_reg, col_reg}==19'b0111001000100000100)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111001000100000101)) color_data = 12'b000000110000;
		if(({row_reg, col_reg}==19'b0111001000100000110)) color_data = 12'b001001000001;
		if(({row_reg, col_reg}==19'b0111001000100000111)) color_data = 12'b010001110100;
		if(({row_reg, col_reg}==19'b0111001000100001000)) color_data = 12'b101011011010;
		if(({row_reg, col_reg}==19'b0111001000100001001)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111001000100001010)) color_data = 12'b100010100111;
		if(({row_reg, col_reg}==19'b0111001000100001011)) color_data = 12'b100110111000;
		if(({row_reg, col_reg}==19'b0111001000100001100)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111001000100001101)) color_data = 12'b010001110100;
		if(({row_reg, col_reg}==19'b0111001000100001110)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0111001000100001111) && ({row_reg, col_reg}<19'b0111001000100011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000100011001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001000100011010)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0111001000100011011)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0111001000100011100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001000100011101)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0111001000100011110)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==19'b0111001000100011111)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0111001000100100000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0111001000100100001)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001000100100010)) color_data = 12'b000101000010;
		if(({row_reg, col_reg}==19'b0111001000100100011)) color_data = 12'b010001100100;
		if(({row_reg, col_reg}==19'b0111001000100100100)) color_data = 12'b001001000010;
		if(({row_reg, col_reg}>=19'b0111001000100100101) && ({row_reg, col_reg}<19'b0111001000100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000100100111)) color_data = 12'b000100110001;
		if(({row_reg, col_reg}==19'b0111001000100101000)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001000100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000100101010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001000100101011)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0111001000100101100)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0111001000100101101)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0111001000100101110)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001000100101111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001000100110000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0111001000100110001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001000100110010) && ({row_reg, col_reg}<19'b0111001000100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000100110100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001000100110101) && ({row_reg, col_reg}<19'b0111001000100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000100110111)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001000100111000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001000100111001)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0111001000100111010)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==19'b0111001000100111011)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==19'b0111001000100111100)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==19'b0111001000100111101)) color_data = 12'b101111011101;
		if(({row_reg, col_reg}==19'b0111001000100111110)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==19'b0111001000100111111)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0111001000101000000)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111001000101000001)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==19'b0111001000101000010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001000101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000101000100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001000101000101)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0111001000101000110)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111001000101000111)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0111001000101001000)) color_data = 12'b011010000110;
		if(({row_reg, col_reg}==19'b0111001000101001001)) color_data = 12'b000000110001;
		if(({row_reg, col_reg}==19'b0111001000101001010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001000101001011)) color_data = 12'b011010000110;
		if(({row_reg, col_reg}==19'b0111001000101001100)) color_data = 12'b101011011011;
		if(({row_reg, col_reg}==19'b0111001000101001101)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111001000101001110)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==19'b0111001000101001111)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0111001000101010000)) color_data = 12'b010101110101;
		if(({row_reg, col_reg}==19'b0111001000101010001)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001000101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000101010011)) color_data = 12'b001001000010;
		if(({row_reg, col_reg}==19'b0111001000101010100)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0111001000101010101)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==19'b0111001000101010110)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0111001000101010111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001000101011000)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0111001000101011001)) color_data = 12'b101011011011;
		if(({row_reg, col_reg}==19'b0111001000101011010)) color_data = 12'b010110000110;
		if(({row_reg, col_reg}==19'b0111001000101011011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001000101011100)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0111001000101011101)) color_data = 12'b100110111001;
		if(({row_reg, col_reg}==19'b0111001000101011110)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==19'b0111001000101011111)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==19'b0111001000101100000)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==19'b0111001000101100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111001000101100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111001000101100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111001000101100100) && ({row_reg, col_reg}<19'b0111001000101100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001000101100110) && ({row_reg, col_reg}<19'b0111001000101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111001000101101000) && ({row_reg, col_reg}<19'b0111001000101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000101110001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111001000101110010) && ({row_reg, col_reg}<19'b0111001000101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001000101111010)) color_data = 12'b010001000000;
		if(({row_reg, col_reg}==19'b0111001000101111011)) color_data = 12'b011001110011;
		if(({row_reg, col_reg}==19'b0111001000101111100)) color_data = 12'b101010110110;
		if(({row_reg, col_reg}==19'b0111001000101111101)) color_data = 12'b110111101001;
		if(({row_reg, col_reg}==19'b0111001000101111110)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}==19'b0111001000101111111)) color_data = 12'b110011011000;
		if(({row_reg, col_reg}==19'b0111001000110000000)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0111001000110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001000110000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111001000110000011) && ({row_reg, col_reg}<19'b0111001001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001001001010001) && ({row_reg, col_reg}<19'b0111001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111001001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111001001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111001010000000000) && ({row_reg, col_reg}<19'b0111001010011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111001010011110011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001010011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010011110101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001010011110110)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0111001010011110111)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==19'b0111001010011111000)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==19'b0111001010011111001)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==19'b0111001010011111010)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==19'b0111001010011111011)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==19'b0111001010011111100)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==19'b0111001010011111101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001010011111110)) color_data = 12'b000001000011;
		if(({row_reg, col_reg}==19'b0111001010011111111)) color_data = 12'b010110010111;
		if(({row_reg, col_reg}==19'b0111001010100000000)) color_data = 12'b100010111000;
		if(({row_reg, col_reg}==19'b0111001010100000001)) color_data = 12'b011010000101;
		if(({row_reg, col_reg}==19'b0111001010100000010)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0111001010100000011)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0111001010100000100) && ({row_reg, col_reg}<19'b0111001010100000110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001010100000110)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001010100000111)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111001010100001000)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}>=19'b0111001010100001001) && ({row_reg, col_reg}<19'b0111001010100001011)) color_data = 12'b001001000001;
		if(({row_reg, col_reg}==19'b0111001010100001011)) color_data = 12'b001001010010;
		if(({row_reg, col_reg}==19'b0111001010100001100)) color_data = 12'b001101010010;
		if(({row_reg, col_reg}==19'b0111001010100001101)) color_data = 12'b000101000001;
		if(({row_reg, col_reg}==19'b0111001010100001110)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0111001010100001111) && ({row_reg, col_reg}<19'b0111001010100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010100011000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111001010100011001) && ({row_reg, col_reg}<19'b0111001010100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010100011110)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0111001010100011111)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==19'b0111001010100100000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001010100100001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001010100100010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001010100100011)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0111001010100100100)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111001010100100101) && ({row_reg, col_reg}<19'b0111001010100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010100100111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001010100101000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111001010100101001) && ({row_reg, col_reg}<19'b0111001010100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010100101011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001010100101100)) color_data = 12'b001001000010;
		if(({row_reg, col_reg}==19'b0111001010100101101)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0111001010100101110) && ({row_reg, col_reg}<19'b0111001010100110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001010100110110) && ({row_reg, col_reg}<19'b0111001010100111000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001010100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010100111001)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}>=19'b0111001010100111010) && ({row_reg, col_reg}<19'b0111001010100111100)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}>=19'b0111001010100111100) && ({row_reg, col_reg}<19'b0111001010100111110)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==19'b0111001010100111110)) color_data = 12'b010001100101;
		if(({row_reg, col_reg}>=19'b0111001010100111111) && ({row_reg, col_reg}<19'b0111001010101000001)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0111001010101000001)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001010101000010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001010101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001010101000100) && ({row_reg, col_reg}<19'b0111001010101001000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001010101001000)) color_data = 12'b001001000010;
		if(({row_reg, col_reg}>=19'b0111001010101001001) && ({row_reg, col_reg}<19'b0111001010101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010101001011)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0111001010101001100)) color_data = 12'b011010010111;
		if(({row_reg, col_reg}==19'b0111001010101001101)) color_data = 12'b100010101000;
		if(({row_reg, col_reg}==19'b0111001010101001110)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0111001010101001111)) color_data = 12'b010001110101;
		if(({row_reg, col_reg}==19'b0111001010101010000)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}==19'b0111001010101010001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001010101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010101010011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001010101010100)) color_data = 12'b010001100100;
		if(({row_reg, col_reg}==19'b0111001010101010101)) color_data = 12'b010101110101;
		if(({row_reg, col_reg}==19'b0111001010101010110)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0111001010101010111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001010101011000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001010101011001)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0111001010101011010)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0111001010101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010101011100)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001010101011101)) color_data = 12'b010001100101;
		if(({row_reg, col_reg}==19'b0111001010101011110)) color_data = 12'b011110010111;
		if(({row_reg, col_reg}==19'b0111001010101011111)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==19'b0111001010101100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001010101100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001010101100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001010101100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111001010101100100) && ({row_reg, col_reg}<19'b0111001010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001010101111000) && ({row_reg, col_reg}<19'b0111001010101111010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001010101111010) && ({row_reg, col_reg}<19'b0111001010101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001010101111100)) color_data = 12'b001101000000;
		if(({row_reg, col_reg}==19'b0111001010101111101)) color_data = 12'b101010110110;
		if(({row_reg, col_reg}==19'b0111001010101111110)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==19'b0111001010101111111)) color_data = 12'b111011111011;
		if(({row_reg, col_reg}==19'b0111001010110000000)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==19'b0111001010110000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111001010110000010) && ({row_reg, col_reg}<19'b0111001010110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001010110000100) && ({row_reg, col_reg}<19'b0111001010110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111001010110000110) && ({row_reg, col_reg}<19'b0111001011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001011001010001) && ({row_reg, col_reg}<19'b0111001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111001011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111001011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111001100000000000) && ({row_reg, col_reg}<19'b0111001100011110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100011110101)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001100011110110)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001100011110111)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0111001100011111000)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==19'b0111001100011111001)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==19'b0111001100011111010)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==19'b0111001100011111011)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==19'b0111001100011111100)) color_data = 12'b001001010100;
		if(({row_reg, col_reg}==19'b0111001100011111101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100011111110)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001100011111111)) color_data = 12'b001001010011;
		if(({row_reg, col_reg}==19'b0111001100100000000)) color_data = 12'b001101010011;
		if(({row_reg, col_reg}==19'b0111001100100000001)) color_data = 12'b001001000010;
		if(({row_reg, col_reg}==19'b0111001100100000010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}>=19'b0111001100100000011) && ({row_reg, col_reg}<19'b0111001100100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001100100000110) && ({row_reg, col_reg}<19'b0111001100100001000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001100100001000) && ({row_reg, col_reg}<19'b0111001100100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100100001100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001100100001101) && ({row_reg, col_reg}<19'b0111001100100001111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001100100001111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001100100010000) && ({row_reg, col_reg}<19'b0111001100100011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100100011000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001100100011001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001100100011010) && ({row_reg, col_reg}<19'b0111001100100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100100011111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100100100000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111001100100100001) && ({row_reg, col_reg}<19'b0111001100100100011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100100100011)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001100100100100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001100100100101) && ({row_reg, col_reg}<19'b0111001100100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100100100111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001100100101000)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0111001100100101001) && ({row_reg, col_reg}<19'b0111001100100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001100100101011) && ({row_reg, col_reg}<19'b0111001100100101101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001100100101101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100100101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100100101111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111001100100110000) && ({row_reg, col_reg}<19'b0111001100100110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100100110010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001100100110011) && ({row_reg, col_reg}<19'b0111001100100111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100100111001)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001100100111010)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0111001100100111011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100100111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100100111101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001100100111110) && ({row_reg, col_reg}<19'b0111001100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001100101000000) && ({row_reg, col_reg}<19'b0111001100101000100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100101000100)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001100101000101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001100101000110) && ({row_reg, col_reg}<19'b0111001100101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100101001000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100101001001)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001100101001010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001100101001011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100101001100)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0111001100101001101)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==19'b0111001100101001110)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0111001100101001111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001100101010000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001100101010001) && ({row_reg, col_reg}<19'b0111001100101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100101010011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100101010100)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0111001100101010101)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0111001100101010110)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111001100101010111) && ({row_reg, col_reg}<19'b0111001100101011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100101011001)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0111001100101011010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100101011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100101011100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001100101011101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001100101011110)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0111001100101011111)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}>=19'b0111001100101100000) && ({row_reg, col_reg}<19'b0111001100101100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111001100101100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111001100101100011) && ({row_reg, col_reg}<19'b0111001100101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001100101111000) && ({row_reg, col_reg}<19'b0111001100101111010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=19'b0111001100101111010) && ({row_reg, col_reg}<19'b0111001100101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100101111101)) color_data = 12'b011101110011;
		if(({row_reg, col_reg}==19'b0111001100101111110)) color_data = 12'b110111101010;
		if(({row_reg, col_reg}==19'b0111001100101111111)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0111001100110000000)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==19'b0111001100110000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111001100110000010) && ({row_reg, col_reg}<19'b0111001100110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001100110000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111001100110000101) && ({row_reg, col_reg}<19'b0111001101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001101001010001) && ({row_reg, col_reg}<19'b0111001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111001101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111001101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111001110000000000) && ({row_reg, col_reg}<19'b0111001110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110011110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111001110011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111001110011110010) && ({row_reg, col_reg}<19'b0111001110011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110011111010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001110011111011) && ({row_reg, col_reg}<19'b0111001110011111101)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111001110011111101) && ({row_reg, col_reg}<19'b0111001110011111111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110011111111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111001110100000000) && ({row_reg, col_reg}<19'b0111001110100000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001110100000011) && ({row_reg, col_reg}<19'b0111001110100000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001110100000101) && ({row_reg, col_reg}<19'b0111001110100000111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001110100001000) && ({row_reg, col_reg}<19'b0111001110100001010)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001110100001010)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001110100001011) && ({row_reg, col_reg}<19'b0111001110100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001110100001101) && ({row_reg, col_reg}<19'b0111001110100001111)) color_data = 12'b000000100000;
		if(({row_reg, col_reg}==19'b0111001110100001111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001110100010000) && ({row_reg, col_reg}<19'b0111001110100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001110100011010) && ({row_reg, col_reg}<19'b0111001110100011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111001110100011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111001110100011101) && ({row_reg, col_reg}<19'b0111001110100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110100011111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110100100000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111001110100100001) && ({row_reg, col_reg}<19'b0111001110100100011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110100100011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001110100100100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110100100110)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110100100111)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0111001110100101000)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0111001110100101001) && ({row_reg, col_reg}<19'b0111001110100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001110100101011) && ({row_reg, col_reg}<19'b0111001110100101101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110100101110)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}==19'b0111001110100101111)) color_data = 12'b001001000011;
		if(({row_reg, col_reg}==19'b0111001110100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110100110001)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001110100110010)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0111001110100110011)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111001110100110100) && ({row_reg, col_reg}<19'b0111001110100111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110100111000)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001110100111001)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0111001110100111010)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111001110100111011) && ({row_reg, col_reg}<19'b0111001110100111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110100111101)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0111001110100111110)) color_data = 12'b001000110010;
		if(({row_reg, col_reg}==19'b0111001110100111111)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}==19'b0111001110101000000)) color_data = 12'b000100100010;
		if(({row_reg, col_reg}==19'b0111001110101000001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001110101000010) && ({row_reg, col_reg}<19'b0111001110101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110101000111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110101001001)) color_data = 12'b001101010100;
		if(({row_reg, col_reg}==19'b0111001110101001010)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==19'b0111001110101001011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110101001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110101001101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110101001110)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}>=19'b0111001110101001111) && ({row_reg, col_reg}<19'b0111001110101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110101010101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111001110101010110) && ({row_reg, col_reg}<19'b0111001110101011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110101011000)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110101011001)) color_data = 12'b000000100001;
		if(({row_reg, col_reg}>=19'b0111001110101011010) && ({row_reg, col_reg}<19'b0111001110101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110101011100)) color_data = 12'b000100110010;
		if(({row_reg, col_reg}>=19'b0111001110101011101) && ({row_reg, col_reg}<19'b0111001110101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110101011111)) color_data = 12'b000100100001;
		if(({row_reg, col_reg}==19'b0111001110101100000)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111001110101100001) && ({row_reg, col_reg}<19'b0111001110101100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111001110101100011) && ({row_reg, col_reg}<19'b0111001110101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001110101100101) && ({row_reg, col_reg}<19'b0111001110101100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111001110101100111) && ({row_reg, col_reg}<19'b0111001110101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110101111001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0111001110101111010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=19'b0111001110101111011) && ({row_reg, col_reg}<19'b0111001110101111101)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111001110101111101)) color_data = 12'b010101100011;
		if(({row_reg, col_reg}==19'b0111001110101111110)) color_data = 12'b110011001001;
		if(({row_reg, col_reg}==19'b0111001110101111111)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==19'b0111001110110000000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=19'b0111001110110000001) && ({row_reg, col_reg}<19'b0111001110110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001110110000011) && ({row_reg, col_reg}<19'b0111001110110000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111001110110000101) && ({row_reg, col_reg}<19'b0111001110110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111001110110000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111001110110001000) && ({row_reg, col_reg}<19'b0111001111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111001111001010001) && ({row_reg, col_reg}<19'b0111001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111001111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111001111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111010000000000000) && ({row_reg, col_reg}<19'b0111010000011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010000011111101) && ({row_reg, col_reg}<19'b0111010000011111111)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111010000011111111) && ({row_reg, col_reg}<19'b0111010000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111010000101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0111010000101111001)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}>=19'b0111010000101111010) && ({row_reg, col_reg}<19'b0111010000101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111010000101111100)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==19'b0111010000101111101)) color_data = 12'b001100110001;
		if(({row_reg, col_reg}==19'b0111010000101111110)) color_data = 12'b010101100011;
		if(({row_reg, col_reg}==19'b0111010000101111111)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=19'b0111010000110000000) && ({row_reg, col_reg}<19'b0111010000110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010000110110110) && ({row_reg, col_reg}<19'b0111010000110111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111010000110111000) && ({row_reg, col_reg}<19'b0111010000110111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111010000110111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111010000111000000) && ({row_reg, col_reg}<19'b0111010001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010001001010001) && ({row_reg, col_reg}<19'b0111010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111010001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111010001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111010010000000000) && ({row_reg, col_reg}<19'b0111010010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111010010101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0111010010101111001) && ({row_reg, col_reg}<19'b0111010010101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111010010101111101)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==19'b0111010010101111110)) color_data = 12'b001000110001;
		if(({row_reg, col_reg}==19'b0111010010101111111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=19'b0111010010110000000) && ({row_reg, col_reg}<19'b0111010011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010011001010001) && ({row_reg, col_reg}<19'b0111010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111010011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111010011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111010100000000000) && ({row_reg, col_reg}<19'b0111010100011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111010100011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0111010100011110010) && ({row_reg, col_reg}<19'b0111010100101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111010100101111000)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=19'b0111010100101111001) && ({row_reg, col_reg}<19'b0111010100110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010100110111000) && ({row_reg, col_reg}<19'b0111010100110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111010100110111100) && ({row_reg, col_reg}<19'b0111010101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010101001010001) && ({row_reg, col_reg}<19'b0111010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111010101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111010101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111010110000000000) && ({row_reg, col_reg}<19'b0111010110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010110011110000) && ({row_reg, col_reg}<19'b0111010110011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0111010110011110100) && ({row_reg, col_reg}<19'b0111010110100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010110100100001) && ({row_reg, col_reg}<19'b0111010110100101111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111010110100101111) && ({row_reg, col_reg}<19'b0111010110101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010110101000001) && ({row_reg, col_reg}<19'b0111010110101011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111010110101011111) && ({row_reg, col_reg}<19'b0111010110110111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111010110110111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111010110110111101) && ({row_reg, col_reg}<19'b0111010111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111010111001010001) && ({row_reg, col_reg}<19'b0111010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111010111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111010111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111011000000000000) && ({row_reg, col_reg}<19'b0111011000011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011000011110000) && ({row_reg, col_reg}<19'b0111011000011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0111011000011110101) && ({row_reg, col_reg}<19'b0111011000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011000100010001) && ({row_reg, col_reg}<19'b0111011000100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0111011000100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011000100100000) && ({row_reg, col_reg}<19'b0111011000100101111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011000100101111) && ({row_reg, col_reg}<19'b0111011000101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011000101000000) && ({row_reg, col_reg}<19'b0111011000101011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011000101011111) && ({row_reg, col_reg}<19'b0111011000101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011000101111011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111011000101111100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111011000101111101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011000101111110) && ({row_reg, col_reg}<19'b0111011000110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011000110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111011000110111110) && ({row_reg, col_reg}<19'b0111011001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011001001010001) && ({row_reg, col_reg}<19'b0111011001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111011001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111011001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111011010000000000) && ({row_reg, col_reg}<19'b0111011010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011010011110000) && ({row_reg, col_reg}<19'b0111011010011110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0111011010011110101) && ({row_reg, col_reg}<19'b0111011010100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011010100010001) && ({row_reg, col_reg}<19'b0111011010100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0111011010100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011010100100000) && ({row_reg, col_reg}<19'b0111011010100110000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011010100110000) && ({row_reg, col_reg}<19'b0111011010101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011010101000000) && ({row_reg, col_reg}<19'b0111011010101100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011010101100000) && ({row_reg, col_reg}<19'b0111011010101111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011010101111010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111011010101111011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111011010101111100) && ({row_reg, col_reg}<19'b0111011010101111111)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0111011010101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111011010110000000) && ({row_reg, col_reg}<19'b0111011010110110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011010110110011) && ({row_reg, col_reg}<19'b0111011010110110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111011010110110110) && ({row_reg, col_reg}<19'b0111011010110111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011010110111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111011010110111001) && ({row_reg, col_reg}<19'b0111011010110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011010110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111011010110111110) && ({row_reg, col_reg}<19'b0111011011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011011001010001) && ({row_reg, col_reg}<19'b0111011011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111011011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111011011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111011100000000000) && ({row_reg, col_reg}<19'b0111011100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011100011110000) && ({row_reg, col_reg}<19'b0111011100011110110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0111011100011110110) && ({row_reg, col_reg}<19'b0111011100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011100100010000) && ({row_reg, col_reg}<19'b0111011100100100000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0111011100100100000) && ({row_reg, col_reg}<19'b0111011100100110000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011100100110000) && ({row_reg, col_reg}<19'b0111011100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011100101000000) && ({row_reg, col_reg}<19'b0111011100101100000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011100101100000) && ({row_reg, col_reg}<19'b0111011100101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011100101111001) && ({row_reg, col_reg}<19'b0111011100101111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111011100101111110)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}==19'b0111011100101111111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111011100110000000) && ({row_reg, col_reg}<19'b0111011100110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011100110110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111011100110110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111011100110110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111011100110110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111011100110110100) && ({row_reg, col_reg}<19'b0111011100110110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111011100110110110) && ({row_reg, col_reg}<19'b0111011100110111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111011100110111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011100110111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111011100110111010) && ({row_reg, col_reg}<19'b0111011100110111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011100110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111011100110111110) && ({row_reg, col_reg}<19'b0111011101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011101001010001) && ({row_reg, col_reg}<19'b0111011101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111011101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111011101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111011110000000000) && ({row_reg, col_reg}<19'b0111011110011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011110011110000) && ({row_reg, col_reg}<19'b0111011110011110100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0111011110011110100) && ({row_reg, col_reg}<19'b0111011110100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011110100010001) && ({row_reg, col_reg}<19'b0111011110100011111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0111011110100011111) && ({row_reg, col_reg}<19'b0111011110100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011110100100001) && ({row_reg, col_reg}<19'b0111011110100101111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011110100101111) && ({row_reg, col_reg}<19'b0111011110101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011110101000001) && ({row_reg, col_reg}<19'b0111011110101011111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011110101011111) && ({row_reg, col_reg}<19'b0111011110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011110101111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111011110101111001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011110101111010) && ({row_reg, col_reg}<19'b0111011110101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011110101111110) && ({row_reg, col_reg}<19'b0111011110110000000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111011110110000000) && ({row_reg, col_reg}<19'b0111011110110110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011110110110000)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==19'b0111011110110110001)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==19'b0111011110110110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==19'b0111011110110110011)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}>=19'b0111011110110110100) && ({row_reg, col_reg}<19'b0111011110110110110)) color_data = 12'b110111001101;
		if(({row_reg, col_reg}==19'b0111011110110110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111011110110110111)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0111011110110111000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==19'b0111011110110111001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==19'b0111011110110111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111011110110111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111011110110111100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111011110110111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111011110110111110) && ({row_reg, col_reg}<19'b0111011111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111011111001010001) && ({row_reg, col_reg}<19'b0111011111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111011111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111011111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111100000000000000) && ({row_reg, col_reg}<19'b0111100000010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100000010101011) && ({row_reg, col_reg}<19'b0111100000010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000010101110) && ({row_reg, col_reg}<19'b0111100000010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000010111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100000010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000010111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100000010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100000010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000010111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111100000010111110) && ({row_reg, col_reg}<19'b0111100000011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100000011000101) && ({row_reg, col_reg}<19'b0111100000011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000011000111) && ({row_reg, col_reg}<19'b0111100000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000011011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100000011011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000011011111) && ({row_reg, col_reg}<19'b0111100000011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000011100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100000011100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100000011100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000011100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100000011100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111100000011100111) && ({row_reg, col_reg}<19'b0111100000011110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000011110001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=19'b0111100000011110010) && ({row_reg, col_reg}<19'b0111100000011110100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==19'b0111100000011110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000011110101) && ({row_reg, col_reg}<19'b0111100000011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100000011111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100000011111001) && ({row_reg, col_reg}<19'b0111100000011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100000011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000011111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100000011111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111100000011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100000100000000) && ({row_reg, col_reg}<19'b0111100000100001000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100000100001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100000100001001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111100000100001010) && ({row_reg, col_reg}<19'b0111100000100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100000100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100000100001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100000100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000100010001) && ({row_reg, col_reg}<19'b0111100000100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000100100001) && ({row_reg, col_reg}<19'b0111100000100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100000100100011) && ({row_reg, col_reg}<19'b0111100000100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000100100101) && ({row_reg, col_reg}<19'b0111100000100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000100100111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0111100000100101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000100101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100000100101010)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}==19'b0111100000100101011)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111100000100101100) && ({row_reg, col_reg}<19'b0111100000100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000100101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100000100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100000100110001) && ({row_reg, col_reg}<19'b0111100000100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100000100110011) && ({row_reg, col_reg}<19'b0111100000100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000100110101) && ({row_reg, col_reg}<19'b0111100000100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000100111000) && ({row_reg, col_reg}<19'b0111100000101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000101000010)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111100000101000011) && ({row_reg, col_reg}<19'b0111100000101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000101000101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100000101000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100000101000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000101001000)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0111100000101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000101001010) && ({row_reg, col_reg}<19'b0111100000101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000101010010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100000101010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100000101010100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111100000101010101) && ({row_reg, col_reg}<19'b0111100000101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000101101001) && ({row_reg, col_reg}<19'b0111100000101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100000101110100) && ({row_reg, col_reg}<19'b0111100000101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000101110110) && ({row_reg, col_reg}<19'b0111100000101111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000101111010) && ({row_reg, col_reg}<19'b0111100000101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000101111100)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==19'b0111100000101111101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100000101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000101111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100000110000000) && ({row_reg, col_reg}<19'b0111100000110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000110010001) && ({row_reg, col_reg}<19'b0111100000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100000110010101) && ({row_reg, col_reg}<19'b0111100000110011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100000110011000) && ({row_reg, col_reg}<19'b0111100000110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000110101000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100000110101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100000110101010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100000110101011)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111100000110101100)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111100000110101101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0111100000110101110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100000110101111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==19'b0111100000110110000)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0111100000110110001)) color_data = 12'b111010111101;
		if(({row_reg, col_reg}==19'b0111100000110110010)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0111100000110110011)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0111100000110110100)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==19'b0111100000110110101)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==19'b0111100000110110110)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==19'b0111100000110110111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==19'b0111100000110111000)) color_data = 12'b110111001101;
		if(({row_reg, col_reg}==19'b0111100000110111001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==19'b0111100000110111010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0111100000110111011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100000110111100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0111100000110111101)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111100000110111110) && ({row_reg, col_reg}<19'b0111100001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100001001010001) && ({row_reg, col_reg}<19'b0111100001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111100001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111100010000000000) && ({row_reg, col_reg}<19'b0111100010010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100010010101011) && ({row_reg, col_reg}<19'b0111100010010101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010010101110) && ({row_reg, col_reg}<19'b0111100010010110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010010110001) && ({row_reg, col_reg}<19'b0111100010010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010010111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010010111010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100010010111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100010010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010010111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100010010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010010111111) && ({row_reg, col_reg}<19'b0111100010011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010011000110) && ({row_reg, col_reg}<19'b0111100010011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010011011001) && ({row_reg, col_reg}<19'b0111100010011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010011011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010011011100) && ({row_reg, col_reg}<19'b0111100010011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010011011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111100010011100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010011100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100010011100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111100010011100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111100010011100100) && ({row_reg, col_reg}<19'b0111100010011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010011100111) && ({row_reg, col_reg}<19'b0111100010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010011110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100010011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010011110010) && ({row_reg, col_reg}<19'b0111100010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010011111001) && ({row_reg, col_reg}<19'b0111100010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010011111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111100010011111111) && ({row_reg, col_reg}<19'b0111100010100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010100001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010100001010) && ({row_reg, col_reg}<19'b0111100010100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100010100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010100001101) && ({row_reg, col_reg}<19'b0111100010100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100010100001111) && ({row_reg, col_reg}<19'b0111100010100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010100010001) && ({row_reg, col_reg}<19'b0111100010100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100010100100011) && ({row_reg, col_reg}<19'b0111100010100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010100100101) && ({row_reg, col_reg}<19'b0111100010100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010100100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100010100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100010100101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100010100101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111100010100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111100010100101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100010100101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100010100101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100010100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100010100110001) && ({row_reg, col_reg}<19'b0111100010100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100010100110011) && ({row_reg, col_reg}<19'b0111100010100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010100110101) && ({row_reg, col_reg}<19'b0111100010101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100010101000010) && ({row_reg, col_reg}<19'b0111100010101000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100010101000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010101000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100010101000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100010101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100010101001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100010101001010) && ({row_reg, col_reg}<19'b0111100010101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010101001101) && ({row_reg, col_reg}<19'b0111100010101001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100010101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010101010000) && ({row_reg, col_reg}<19'b0111100010101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010101101010) && ({row_reg, col_reg}<19'b0111100010101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100010101101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010101101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100010101101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010101110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100010101110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100010101110010) && ({row_reg, col_reg}<19'b0111100010101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010101111101) && ({row_reg, col_reg}<19'b0111100010101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010101111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100010110000000) && ({row_reg, col_reg}<19'b0111100010110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100010110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100010110011000) && ({row_reg, col_reg}<19'b0111100010110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100010110100001) && ({row_reg, col_reg}<19'b0111100010110101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100010110101000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0111100010110101001) && ({row_reg, col_reg}<19'b0111100010110101011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100010110101011)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111100010110101100)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111100010110101101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100010110101110)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111100010110101111)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==19'b0111100010110110000)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==19'b0111100010110110001)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}==19'b0111100010110110010)) color_data = 12'b100001010111;
		if(({row_reg, col_reg}==19'b0111100010110110011)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==19'b0111100010110110100)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0111100010110110101)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==19'b0111100010110110110)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111100010110110111)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0111100010110111000)) color_data = 12'b110111001101;
		if(({row_reg, col_reg}==19'b0111100010110111001)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==19'b0111100010110111010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0111100010110111011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100010110111100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0111100010110111101) && ({row_reg, col_reg}<19'b0111100010110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111100010110111111) && ({row_reg, col_reg}<19'b0111100011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100011001010001) && ({row_reg, col_reg}<19'b0111100011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111100011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111100100000000000) && ({row_reg, col_reg}<19'b0111100100010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100100010110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100100010111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100010111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100100010111011) && ({row_reg, col_reg}<19'b0111100100010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100100010111110) && ({row_reg, col_reg}<19'b0111100100011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100100011000010) && ({row_reg, col_reg}<19'b0111100100011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100011000101) && ({row_reg, col_reg}<19'b0111100100011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100100011011001) && ({row_reg, col_reg}<19'b0111100100011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100011011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100100011011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100011011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100100011011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100100011100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100100011100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100100011100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100100011100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111100100011100100) && ({row_reg, col_reg}<19'b0111100100011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100011100111) && ({row_reg, col_reg}<19'b0111100100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100011110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100100011110001) && ({row_reg, col_reg}<19'b0111100100011110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100011110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100100011110101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100100011110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100100011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100100011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100100011111010) && ({row_reg, col_reg}<19'b0111100100011111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111100100011111100) && ({row_reg, col_reg}<19'b0111100100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100011111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100100011111111) && ({row_reg, col_reg}<19'b0111100100100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100100100001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100100100001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100100100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100100100001101) && ({row_reg, col_reg}<19'b0111100100100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100100001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100100100010000) && ({row_reg, col_reg}<19'b0111100100100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100100100100011) && ({row_reg, col_reg}<19'b0111100100100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100100100101) && ({row_reg, col_reg}<19'b0111100100100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100100100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100100100101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111100100100101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111100100100101010) && ({row_reg, col_reg}<19'b0111100100100101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100100100101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100100100101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100100100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100100100110001) && ({row_reg, col_reg}<19'b0111100100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100100100110011) && ({row_reg, col_reg}<19'b0111100100100110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100100110101) && ({row_reg, col_reg}<19'b0111100100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100101000001) && ({row_reg, col_reg}<19'b0111100100101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100101000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100100101000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111100100101000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111100100101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100100101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111100100101001000) && ({row_reg, col_reg}<19'b0111100100101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100100101001011) && ({row_reg, col_reg}<19'b0111100100101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100101001101) && ({row_reg, col_reg}<19'b0111100100101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100101010001) && ({row_reg, col_reg}<19'b0111100100101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100101011000) && ({row_reg, col_reg}<19'b0111100100101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100101101010) && ({row_reg, col_reg}<19'b0111100100101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100101101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111100100101101101) && ({row_reg, col_reg}<19'b0111100100101101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100100101101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111100100101110000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100100101110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100100101110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111100100101110011) && ({row_reg, col_reg}<19'b0111100100101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100100101111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100100101111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100100101111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100101111011) && ({row_reg, col_reg}<19'b0111100100101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100100101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100110000000) && ({row_reg, col_reg}<19'b0111100100110010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100100110010001) && ({row_reg, col_reg}<19'b0111100100110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100100110010100) && ({row_reg, col_reg}<19'b0111100100110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100100110100001) && ({row_reg, col_reg}<19'b0111100100110101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100100110101000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0111100100110101001) && ({row_reg, col_reg}<19'b0111100100110101011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100100110101011)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111100100110101100)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111100100110101101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100100110101110)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111100100110101111)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}>=19'b0111100100110110000) && ({row_reg, col_reg}<19'b0111100100110110010)) color_data = 12'b101110001010;
		if(({row_reg, col_reg}==19'b0111100100110110010)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}>=19'b0111100100110110011) && ({row_reg, col_reg}<19'b0111100100110110110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100100110110110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111100100110110111)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0111100100110111000)) color_data = 12'b110010111101;
		if(({row_reg, col_reg}==19'b0111100100110111001)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==19'b0111100100110111010)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0111100100110111011)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100100110111100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0111100100110111101) && ({row_reg, col_reg}<19'b0111100100110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111100100110111111) && ({row_reg, col_reg}<19'b0111100101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100101001010001) && ({row_reg, col_reg}<19'b0111100101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111100101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111100110000000000) && ({row_reg, col_reg}<19'b0111100110010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110010101001) && ({row_reg, col_reg}<19'b0111100110010110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100110010110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100110010110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100110010110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111100110010110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100110010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100110010110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100110010111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111100110010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110010111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111100110010111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100110010111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110010111110) && ({row_reg, col_reg}<19'b0111100110011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100110011000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100110011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110011000101) && ({row_reg, col_reg}<19'b0111100110011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100110011001000) && ({row_reg, col_reg}<19'b0111100110011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100110011011001) && ({row_reg, col_reg}<19'b0111100110011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100110011011011) && ({row_reg, col_reg}<19'b0111100110011011110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100110011011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100110011011111) && ({row_reg, col_reg}<19'b0111100110011100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110011100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111100110011100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110011100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111100110011100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100110011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110011100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100110011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110011101000) && ({row_reg, col_reg}<19'b0111100110011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110011110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111100110011110100) && ({row_reg, col_reg}<19'b0111100110011110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100110011110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111100110011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100110011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100110011111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100110011111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100110011111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100110011111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100110011111110) && ({row_reg, col_reg}<19'b0111100110100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110100000001) && ({row_reg, col_reg}<19'b0111100110100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100110100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110100001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100110100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110100001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111100110100001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111100110100001101) && ({row_reg, col_reg}<19'b0111100110100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110100010000) && ({row_reg, col_reg}<19'b0111100110100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110100010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110100010011) && ({row_reg, col_reg}<19'b0111100110100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110100100100) && ({row_reg, col_reg}<19'b0111100110100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110100100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100110100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100110100101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111100110100101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100110100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111100110100101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100110100101101) && ({row_reg, col_reg}<19'b0111100110100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110100101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111100110100110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111100110100110001) && ({row_reg, col_reg}<19'b0111100110100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110100110101) && ({row_reg, col_reg}<19'b0111100110101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100110101000001) && ({row_reg, col_reg}<19'b0111100110101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110101000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111100110101000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111100110101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110101000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111100110101001000) && ({row_reg, col_reg}<19'b0111100110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110101010000) && ({row_reg, col_reg}<19'b0111100110101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100110101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111100110101101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100110101101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111100110101101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110101101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111100110101101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100110101110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110101110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111100110101110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100110101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100110101110100) && ({row_reg, col_reg}<19'b0111100110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110101111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100110101111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100110101111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111100110101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110101111101) && ({row_reg, col_reg}<19'b0111100110101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111100110110000000) && ({row_reg, col_reg}<19'b0111100110110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111100110110010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111100110110010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111100110110010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111100110110010111) && ({row_reg, col_reg}<19'b0111100110110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100110110100001) && ({row_reg, col_reg}<19'b0111100110110101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111100110110101000) && ({row_reg, col_reg}<19'b0111100110110101011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111100110110101011) && ({row_reg, col_reg}<19'b0111100110110101101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111100110110101101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100110110101110)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111100110110101111)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==19'b0111100110110110000)) color_data = 12'b110110101100;
		if(({row_reg, col_reg}==19'b0111100110110110001)) color_data = 12'b101110001010;
		if(({row_reg, col_reg}==19'b0111100110110110010)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}>=19'b0111100110110110011) && ({row_reg, col_reg}<19'b0111100110110110110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111100110110110110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111100110110110111)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0111100110110111000)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==19'b0111100110110111001)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}>=19'b0111100110110111010) && ({row_reg, col_reg}<19'b0111100110110111100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100110110111100)) color_data = 12'b000000000010;
		if(({row_reg, col_reg}>=19'b0111100110110111101) && ({row_reg, col_reg}<19'b0111100110110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111100110110111111) && ({row_reg, col_reg}<19'b0111100111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111100111001010001) && ({row_reg, col_reg}<19'b0111100111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111100111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111100111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111101000000000000) && ({row_reg, col_reg}<19'b0111101000010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101000010101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101000010101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111101000010101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000010110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101000010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101000010110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101000010110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111101000010110100) && ({row_reg, col_reg}<19'b0111101000010111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000010111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101000010111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101000010111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101000010111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101000010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101000010111101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101000010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000010111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000011000000) && ({row_reg, col_reg}<19'b0111101000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101000011000011) && ({row_reg, col_reg}<19'b0111101000011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000011000101) && ({row_reg, col_reg}<19'b0111101000011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101000011001000) && ({row_reg, col_reg}<19'b0111101000011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000011011010) && ({row_reg, col_reg}<19'b0111101000011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000011011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101000011011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101000011011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101000011011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101000011100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101000011100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111101000011100010) && ({row_reg, col_reg}<19'b0111101000011100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000011100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111101000011100101) && ({row_reg, col_reg}<19'b0111101000011100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101000011100111) && ({row_reg, col_reg}<19'b0111101000011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000011110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111101000011110100) && ({row_reg, col_reg}<19'b0111101000011110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101000011110110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111101000011110111) && ({row_reg, col_reg}<19'b0111101000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101000011111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101000011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000011111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111101000011111101) && ({row_reg, col_reg}<19'b0111101000011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000011111111) && ({row_reg, col_reg}<19'b0111101000100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101000100001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101000100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000100001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111101000100001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111101000100001101) && ({row_reg, col_reg}<19'b0111101000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000100010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101000100010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101000100010011) && ({row_reg, col_reg}<19'b0111101000100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000100100100) && ({row_reg, col_reg}<19'b0111101000100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000100100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101000100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000100101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101000100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111101000100101011) && ({row_reg, col_reg}<19'b0111101000100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000100101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101000100101110) && ({row_reg, col_reg}<19'b0111101000100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000100110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000100110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101000100110010) && ({row_reg, col_reg}<19'b0111101000100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000100110101) && ({row_reg, col_reg}<19'b0111101000101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000101000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101000101000001) && ({row_reg, col_reg}<19'b0111101000101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000101000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111101000101000101) && ({row_reg, col_reg}<19'b0111101000101000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101000101000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101000101001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101000101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101000101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000101001100) && ({row_reg, col_reg}<19'b0111101000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000101001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111101000101010000) && ({row_reg, col_reg}<19'b0111101000101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101000101010100) && ({row_reg, col_reg}<19'b0111101000101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000101010110) && ({row_reg, col_reg}<19'b0111101000101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101000101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000101101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111101000101101011) && ({row_reg, col_reg}<19'b0111101000101101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000101101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101000101101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101000101101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101000101110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101000101110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101000101110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000101110011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101000101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000101110101) && ({row_reg, col_reg}<19'b0111101000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101000101111000) && ({row_reg, col_reg}<19'b0111101000101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000101111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111101000101111011) && ({row_reg, col_reg}<19'b0111101000101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101000101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000110000000) && ({row_reg, col_reg}<19'b0111101000110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101000110010001) && ({row_reg, col_reg}<19'b0111101000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101000110010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111101000110010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101000110010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111101000110010111) && ({row_reg, col_reg}<19'b0111101000110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101000110100001) && ({row_reg, col_reg}<19'b0111101000110101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111101000110101001) && ({row_reg, col_reg}<19'b0111101000110101011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111101000110101011)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111101000110101100)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111101000110101101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111101000110101110)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111101000110101111)) color_data = 12'b011000110101;
		if(({row_reg, col_reg}==19'b0111101000110110000)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}==19'b0111101000110110001)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==19'b0111101000110110010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111101000110110011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111101000110110100)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111101000110110101)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111101000110110110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0111101000110110111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==19'b0111101000110111000)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==19'b0111101000110111001)) color_data = 12'b010101000110;
		if(({row_reg, col_reg}>=19'b0111101000110111010) && ({row_reg, col_reg}<19'b0111101000110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111101000110111111) && ({row_reg, col_reg}<19'b0111101001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101001001010001) && ({row_reg, col_reg}<19'b0111101001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111101001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111101001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111101010000000000) && ({row_reg, col_reg}<19'b0111101010010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010010101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101010010101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101010010101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111101010010101111) && ({row_reg, col_reg}<19'b0111101010010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010010110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101010010110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101010010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101010010110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101010010111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111101010010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111101010010111010) && ({row_reg, col_reg}<19'b0111101010010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111101010010111101) && ({row_reg, col_reg}<19'b0111101010010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010010111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101010011000000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111101010011000001) && ({row_reg, col_reg}<19'b0111101010011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010011000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010011000101) && ({row_reg, col_reg}<19'b0111101010011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101010011001000) && ({row_reg, col_reg}<19'b0111101010011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010011011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101010011011010) && ({row_reg, col_reg}<19'b0111101010011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010011011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111101010011011101) && ({row_reg, col_reg}<19'b0111101010011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010011011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111101010011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010011100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101010011100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101010011100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101010011100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101010011100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101010011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010011100111) && ({row_reg, col_reg}<19'b0111101010011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010011110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101010011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101010011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101010011110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101010011110101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101010011110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101010011110111) && ({row_reg, col_reg}<19'b0111101010011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101010011111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101010011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010011111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111101010011111101) && ({row_reg, col_reg}<19'b0111101010100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101010100000011) && ({row_reg, col_reg}<19'b0111101010100000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010100000101) && ({row_reg, col_reg}<19'b0111101010100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101010100001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101010100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010100001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101010100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101010100001101) && ({row_reg, col_reg}<19'b0111101010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101010100010001) && ({row_reg, col_reg}<19'b0111101010100010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111101010100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010100010100) && ({row_reg, col_reg}<19'b0111101010100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010100010111) && ({row_reg, col_reg}<19'b0111101010100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010100100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101010100100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101010100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010100101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101010100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010100101011) && ({row_reg, col_reg}<19'b0111101010100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101010100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101010100101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101010100110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101010100110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111101010100110010) && ({row_reg, col_reg}<19'b0111101010101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010101000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111101010101000101) && ({row_reg, col_reg}<19'b0111101010101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010101000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101010101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010101001001) && ({row_reg, col_reg}<19'b0111101010101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010101001100) && ({row_reg, col_reg}<19'b0111101010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010101001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101010101010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101010101010001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010101010010) && ({row_reg, col_reg}<19'b0111101010101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101010101010100) && ({row_reg, col_reg}<19'b0111101010101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010101010110) && ({row_reg, col_reg}<19'b0111101010101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010101101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101010101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101010101101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101010101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010101101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101010101101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111101010101101110) && ({row_reg, col_reg}<19'b0111101010101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010101110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101010101110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101010101110010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101010101110011) && ({row_reg, col_reg}<19'b0111101010101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010101110110) && ({row_reg, col_reg}<19'b0111101010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010101111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111101010101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101010101111011) && ({row_reg, col_reg}<19'b0111101010101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101010101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010101111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010110000000) && ({row_reg, col_reg}<19'b0111101010110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101010110010001) && ({row_reg, col_reg}<19'b0111101010110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101010110010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101010110010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010110010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111101010110010111) && ({row_reg, col_reg}<19'b0111101010110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101010110100001) && ({row_reg, col_reg}<19'b0111101010110101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111101010110101001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111101010110101010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==19'b0111101010110101011)) color_data = 12'b011000110101;
		if(({row_reg, col_reg}==19'b0111101010110101100)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==19'b0111101010110101101)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==19'b0111101010110101110)) color_data = 12'b011000110101;
		if(({row_reg, col_reg}==19'b0111101010110101111)) color_data = 12'b100001010111;
		if(({row_reg, col_reg}==19'b0111101010110110000)) color_data = 12'b101110001010;
		if(({row_reg, col_reg}==19'b0111101010110110001)) color_data = 12'b100001010111;
		if(({row_reg, col_reg}==19'b0111101010110110010)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111101010110110011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111101010110110100)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=19'b0111101010110110101) && ({row_reg, col_reg}<19'b0111101010110110111)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111101010110110111)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0111101010110111000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==19'b0111101010110111001)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}>=19'b0111101010110111010) && ({row_reg, col_reg}<19'b0111101010110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111101010110111111) && ({row_reg, col_reg}<19'b0111101011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101011001010001) && ({row_reg, col_reg}<19'b0111101011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111101011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111101011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111101100000000000) && ({row_reg, col_reg}<19'b0111101100010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100010101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101100010101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101100010101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101100010101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0111101100010110000) && ({row_reg, col_reg}<19'b0111101100010110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101100010110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101100010110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100010110100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101100010110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101100010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100010110111) && ({row_reg, col_reg}<19'b0111101100010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100010111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100010111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101100010111100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101100010111101) && ({row_reg, col_reg}<19'b0111101100010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100010111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101100011000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101100011000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111101100011000010) && ({row_reg, col_reg}<19'b0111101100011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101100011000101) && ({row_reg, col_reg}<19'b0111101100011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100011001000) && ({row_reg, col_reg}<19'b0111101100011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100011011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101100011011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101100011011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100011011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101100011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100011100000) && ({row_reg, col_reg}<19'b0111101100011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100011100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101100011100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101100011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101100011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100011100111) && ({row_reg, col_reg}<19'b0111101100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100011110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101100011110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100011110010) && ({row_reg, col_reg}<19'b0111101100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100011111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101100011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100011111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111101100011111101) && ({row_reg, col_reg}<19'b0111101100100000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100100000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101100100000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111101100100000011) && ({row_reg, col_reg}<19'b0111101100100000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101100100000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111101100100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100100000111) && ({row_reg, col_reg}<19'b0111101100100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100100001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101100100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100100001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101100100001100) && ({row_reg, col_reg}<19'b0111101100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100100001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101100100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111101100100010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101100100010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101100100010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101100100010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111101100100010100) && ({row_reg, col_reg}<19'b0111101100100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100100010111) && ({row_reg, col_reg}<19'b0111101100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101100100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101100100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100100101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101100100101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101100100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101100100101011) && ({row_reg, col_reg}<19'b0111101100100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101100100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100100101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101100100101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101100100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100100110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101100100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100100110011) && ({row_reg, col_reg}<19'b0111101100101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100101000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101100101000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101100101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100101000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111101100101000101) && ({row_reg, col_reg}<19'b0111101100101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100101000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111101100101001000) && ({row_reg, col_reg}<19'b0111101100101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100101001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101100101001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111101100101001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101100101001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101100101001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101100101001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101100101010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100101010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101100101010011) && ({row_reg, col_reg}<19'b0111101100101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100101010110) && ({row_reg, col_reg}<19'b0111101100101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100101101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101100101101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100101101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111101100101101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111101100101101101) && ({row_reg, col_reg}<19'b0111101100101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101100101110100) && ({row_reg, col_reg}<19'b0111101100101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100101110110) && ({row_reg, col_reg}<19'b0111101100101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100101111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101100101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101100101111011) && ({row_reg, col_reg}<19'b0111101100101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100101111110) && ({row_reg, col_reg}<19'b0111101100110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101100110010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101100110010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101100110010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100110010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101100110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101100110011000) && ({row_reg, col_reg}<19'b0111101100110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101100110100001) && ({row_reg, col_reg}<19'b0111101100110101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111101100110101001)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111101100110101010)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==19'b0111101100110101011)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==19'b0111101100110101100)) color_data = 12'b101110001010;
		if(({row_reg, col_reg}>=19'b0111101100110101101) && ({row_reg, col_reg}<19'b0111101100110101111)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==19'b0111101100110101111)) color_data = 12'b101110001010;
		if(({row_reg, col_reg}==19'b0111101100110110000)) color_data = 12'b110010001011;
		if(({row_reg, col_reg}==19'b0111101100110110001)) color_data = 12'b011101000110;
		if(({row_reg, col_reg}>=19'b0111101100110110010) && ({row_reg, col_reg}<19'b0111101100110110100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111101100110110100)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0111101100110110101)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111101100110110110)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111101100110110111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==19'b0111101100110111000)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}==19'b0111101100110111001)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}>=19'b0111101100110111010) && ({row_reg, col_reg}<19'b0111101100110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111101100110111111) && ({row_reg, col_reg}<19'b0111101101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101101001010001) && ({row_reg, col_reg}<19'b0111101101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111101101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111101101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111101110000000000) && ({row_reg, col_reg}<19'b0111101110010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110010101001) && ({row_reg, col_reg}<19'b0111101110010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101110010101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101110010101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101110010101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111101110010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101110010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101110010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110010110011) && ({row_reg, col_reg}<19'b0111101110010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101110010111010) && ({row_reg, col_reg}<19'b0111101110010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101110010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110010111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111101110010111111) && ({row_reg, col_reg}<19'b0111101110011000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110011000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101110011000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101110011000101) && ({row_reg, col_reg}<19'b0111101110011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110011011001) && ({row_reg, col_reg}<19'b0111101110011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110011011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110011011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101110011011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101110011011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111101110011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110011100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101110011100001) && ({row_reg, col_reg}<19'b0111101110011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110011100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110011100100) && ({row_reg, col_reg}<19'b0111101110011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110011100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101110011100111) && ({row_reg, col_reg}<19'b0111101110011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101110011110010) && ({row_reg, col_reg}<19'b0111101110011110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110011110100) && ({row_reg, col_reg}<19'b0111101110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101110011111000) && ({row_reg, col_reg}<19'b0111101110011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101110011111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101110011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110011111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110011111101) && ({row_reg, col_reg}<19'b0111101110011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101110100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110100000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111101110100000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111101110100000011) && ({row_reg, col_reg}<19'b0111101110100000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110100000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101110100000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111101110100000111) && ({row_reg, col_reg}<19'b0111101110100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110100001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101110100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110100001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101110100001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101110100001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101110100001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111101110100010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111101110100010001) && ({row_reg, col_reg}<19'b0111101110100010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110100010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111101110100010100) && ({row_reg, col_reg}<19'b0111101110100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110100010111) && ({row_reg, col_reg}<19'b0111101110100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110100100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110100100001) && ({row_reg, col_reg}<19'b0111101110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110100100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101110100100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101110100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110100101001) && ({row_reg, col_reg}<19'b0111101110100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101110100101011) && ({row_reg, col_reg}<19'b0111101110100101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111101110100101101) && ({row_reg, col_reg}<19'b0111101110100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110100101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101110100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110100110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101110100110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110100110011) && ({row_reg, col_reg}<19'b0111101110100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110100111000) && ({row_reg, col_reg}<19'b0111101110101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101110101000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101110101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101110101000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111101110101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110101000111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101110101001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111101110101001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101110101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110101001011) && ({row_reg, col_reg}<19'b0111101110101001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111101110101001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101110101001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111101110101001111) && ({row_reg, col_reg}<19'b0111101110101010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110101010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101110101010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111101110101010011) && ({row_reg, col_reg}<19'b0111101110101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110101101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111101110101101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110101101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110101101100) && ({row_reg, col_reg}<19'b0111101110101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110101101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111101110101101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111101110101110000) && ({row_reg, col_reg}<19'b0111101110101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110101110010) && ({row_reg, col_reg}<19'b0111101110101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101110101110100) && ({row_reg, col_reg}<19'b0111101110101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110101110110) && ({row_reg, col_reg}<19'b0111101110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110101111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111101110101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111101110101111011) && ({row_reg, col_reg}<19'b0111101110101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110101111110) && ({row_reg, col_reg}<19'b0111101110110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111101110110010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111101110110010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101110110010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110110010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101110110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111101110110011000) && ({row_reg, col_reg}<19'b0111101110110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101110110100001) && ({row_reg, col_reg}<19'b0111101110110101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111101110110101000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111101110110101001)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111101110110101010)) color_data = 12'b100001010111;
		if(({row_reg, col_reg}==19'b0111101110110101011)) color_data = 12'b110110101100;
		if(({row_reg, col_reg}==19'b0111101110110101100)) color_data = 12'b111010111101;
		if(({row_reg, col_reg}>=19'b0111101110110101101) && ({row_reg, col_reg}<19'b0111101110110101111)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}>=19'b0111101110110101111) && ({row_reg, col_reg}<19'b0111101110110110001)) color_data = 12'b110110101100;
		if(({row_reg, col_reg}==19'b0111101110110110001)) color_data = 12'b100001010111;
		if(({row_reg, col_reg}>=19'b0111101110110110010) && ({row_reg, col_reg}<19'b0111101110110110100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111101110110110100)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==19'b0111101110110110101)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==19'b0111101110110110110)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==19'b0111101110110110111)) color_data = 12'b111011001110;
		if(({row_reg, col_reg}==19'b0111101110110111000)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}==19'b0111101110110111001)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}>=19'b0111101110110111010) && ({row_reg, col_reg}<19'b0111101110110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111101110110111111) && ({row_reg, col_reg}<19'b0111101111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111101111001010001) && ({row_reg, col_reg}<19'b0111101111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111101111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111101111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111110000000000000) && ({row_reg, col_reg}<19'b0111110000010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110000010101010) && ({row_reg, col_reg}<19'b0111110000010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111110000010101110) && ({row_reg, col_reg}<19'b0111110000010110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110000010110001) && ({row_reg, col_reg}<19'b0111110000010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000010110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110000010110100) && ({row_reg, col_reg}<19'b0111110000010110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110000010110110) && ({row_reg, col_reg}<19'b0111110000010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110000010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110000010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111110000010111101) && ({row_reg, col_reg}<19'b0111110000010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000010111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000011000000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110000011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000011000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110000011000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000011000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000011001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110000011001010) && ({row_reg, col_reg}<19'b0111110000011001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110000011001100) && ({row_reg, col_reg}<19'b0111110000011011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000011011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111110000011011100) && ({row_reg, col_reg}<19'b0111110000011011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000011011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110000011011111) && ({row_reg, col_reg}<19'b0111110000011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000011100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000011100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110000011100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000011101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110000011101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000011101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000011101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110000011101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110000011101101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110000011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000011110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110000011110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110000011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000011110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110000011110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110000011110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110000011110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110000011110111) && ({row_reg, col_reg}<19'b0111110000011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000011111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110000011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000011111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110000011111101) && ({row_reg, col_reg}<19'b0111110000100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000100000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110000100000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110000100000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111110000100000100) && ({row_reg, col_reg}<19'b0111110000100000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000100000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111110000100000111) && ({row_reg, col_reg}<19'b0111110000100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110000100001001) && ({row_reg, col_reg}<19'b0111110000100001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000100001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110000100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000100001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000100001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110000100001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000100010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110000100010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110000100010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000100010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110000100010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110000100010101) && ({row_reg, col_reg}<19'b0111110000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000100100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110000100100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110000100101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110000100101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110000100101011) && ({row_reg, col_reg}<19'b0111110000100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000100101101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000100101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000100101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110000100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000100110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110000100110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110000100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110000100110110) && ({row_reg, col_reg}<19'b0111110000101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000101000100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000101000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110000101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000101000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110000101001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000101001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110000101001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110000101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000101001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000101001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110000101001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000101010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110000101010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000101010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110000101010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111110000101010100) && ({row_reg, col_reg}<19'b0111110000101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110000101010111) && ({row_reg, col_reg}<19'b0111110000101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110000101101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110000101101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000101101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110000101101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111110000101101101) && ({row_reg, col_reg}<19'b0111110000101101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000101101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110000101110001) && ({row_reg, col_reg}<19'b0111110000101110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110000101110011) && ({row_reg, col_reg}<19'b0111110000101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000101111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110000101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000101111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110000101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000101111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110000101111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110000110000000) && ({row_reg, col_reg}<19'b0111110000110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000110000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110000110000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111110000110000100) && ({row_reg, col_reg}<19'b0111110000110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000110000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000110001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000110001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110000110001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000110001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000110001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110000110001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110000110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000110010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111110000110010010) && ({row_reg, col_reg}<19'b0111110000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110000110010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000110010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110000110010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110000110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110000110011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110000110011001) && ({row_reg, col_reg}<19'b0111110000110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110000110100001) && ({row_reg, col_reg}<19'b0111110000110101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111110000110101000)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0111110000110101001)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==19'b0111110000110101010)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0111110000110101011)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0111110000110101100)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==19'b0111110000110101101)) color_data = 12'b110010011100;
		if(({row_reg, col_reg}==19'b0111110000110101110)) color_data = 12'b111010111101;
		if(({row_reg, col_reg}==19'b0111110000110101111)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}==19'b0111110000110110000)) color_data = 12'b100001010111;
		if(({row_reg, col_reg}==19'b0111110000110110001)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111110000110110010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111110000110110011)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==19'b0111110000110110100)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0111110000110110101)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0111110000110110110)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0111110000110110111)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0111110000110111000)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==19'b0111110000110111001)) color_data = 12'b010101000110;
		if(({row_reg, col_reg}>=19'b0111110000110111010) && ({row_reg, col_reg}<19'b0111110000110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111110000110111111) && ({row_reg, col_reg}<19'b0111110001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110001001010001) && ({row_reg, col_reg}<19'b0111110001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111110001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111110001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111110010000000000) && ({row_reg, col_reg}<19'b0111110010010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110010010101010) && ({row_reg, col_reg}<19'b0111110010010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110010010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111110010010101110) && ({row_reg, col_reg}<19'b0111110010010110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110010010110001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110010010110010) && ({row_reg, col_reg}<19'b0111110010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110010010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110010010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110010010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110010010111111) && ({row_reg, col_reg}<19'b0111110010011000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110010011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010011000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110010011000011) && ({row_reg, col_reg}<19'b0111110010011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010011000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111110010011000110) && ({row_reg, col_reg}<19'b0111110010011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110010011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110010011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110010011011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111110010011011101) && ({row_reg, col_reg}<19'b0111110010011100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010011100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110010011100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110010011100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110010011100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110010011100100) && ({row_reg, col_reg}<19'b0111110010011100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010011100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010011100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110010011101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110010011101010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110010011101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111110010011101100) && ({row_reg, col_reg}<19'b0111110010011101110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110010011101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110010011101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111110010011110000) && ({row_reg, col_reg}<19'b0111110010011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110010011110011) && ({row_reg, col_reg}<19'b0111110010011110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110010011110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111110010011110110) && ({row_reg, col_reg}<19'b0111110010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010011111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110010011111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110010011111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010011111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110010011111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110010011111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110010100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010100000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010100000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110010100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010100000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110010100000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110010100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110010100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010100001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110010100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010100001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010100001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110010100001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111110010100001110) && ({row_reg, col_reg}<19'b0111110010100010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110010100010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110010100010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110010100010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110010100010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010100010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110010100010101) && ({row_reg, col_reg}<19'b0111110010100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110010100100011) && ({row_reg, col_reg}<19'b0111110010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010100100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111110010100101000) && ({row_reg, col_reg}<19'b0111110010100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110010100110000) && ({row_reg, col_reg}<19'b0111110010100110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010100110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110010100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110010100110100) && ({row_reg, col_reg}<19'b0111110010100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110010100110110) && ({row_reg, col_reg}<19'b0111110010101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010101000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110010101000010) && ({row_reg, col_reg}<19'b0111110010101000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110010101000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010101000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110010101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010101000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110010101001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010101001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110010101001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110010101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010101001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110010101001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110010101001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010101010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111110010101010001) && ({row_reg, col_reg}<19'b0111110010101010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110010101010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110010101010101) && ({row_reg, col_reg}<19'b0111110010101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010101101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110010101101010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110010101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010101101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110010101101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010101101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111110010101101111) && ({row_reg, col_reg}<19'b0111110010101110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110010101110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010101110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110010101110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111110010101110110) && ({row_reg, col_reg}<19'b0111110010101111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110010101111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111110010101111001) && ({row_reg, col_reg}<19'b0111110010101111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010101111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110010101111100) && ({row_reg, col_reg}<19'b0111110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010101111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110010101111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110010110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010110000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111110010110000010) && ({row_reg, col_reg}<19'b0111110010110000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0111110010110000100) && ({row_reg, col_reg}<19'b0111110010110000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110010110000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110010110001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110010110001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110010110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010110001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110010110001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110010110001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111110010110001110) && ({row_reg, col_reg}<19'b0111110010110010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010110010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110010110010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110010110010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010110010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110010110010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010110011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110010110011001) && ({row_reg, col_reg}<19'b0111110010110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110010110011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110010110011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110010110011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111110010110011110) && ({row_reg, col_reg}<19'b0111110010110100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110010110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110010110100001) && ({row_reg, col_reg}<19'b0111110010110101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111110010110101000)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111110010110101001)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==19'b0111110010110101010)) color_data = 12'b111011001101;
		if(({row_reg, col_reg}==19'b0111110010110101011)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0111110010110101100)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}>=19'b0111110010110101101) && ({row_reg, col_reg}<19'b0111110010110101111)) color_data = 12'b111010111101;
		if(({row_reg, col_reg}==19'b0111110010110101111)) color_data = 12'b101110001010;
		if(({row_reg, col_reg}==19'b0111110010110110000)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}>=19'b0111110010110110001) && ({row_reg, col_reg}<19'b0111110010110110011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111110010110110011)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==19'b0111110010110110100)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0111110010110110101)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0111110010110110110)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0111110010110110111)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==19'b0111110010110111000)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0111110010110111001)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}>=19'b0111110010110111010) && ({row_reg, col_reg}<19'b0111110010110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111110010110111111) && ({row_reg, col_reg}<19'b0111110011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110011001010001) && ({row_reg, col_reg}<19'b0111110011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111110011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111110011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111110100000000000) && ({row_reg, col_reg}<19'b0111110100010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110100010101010) && ({row_reg, col_reg}<19'b0111110100010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110100010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111110100010101110) && ({row_reg, col_reg}<19'b0111110100010110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0111110100010110000) && ({row_reg, col_reg}<19'b0111110100010110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100010110011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110100010110100) && ({row_reg, col_reg}<19'b0111110100010110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110100010110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110100010110111) && ({row_reg, col_reg}<19'b0111110100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110100010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110100010111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110100010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110100010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100010111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110100010111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100011000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110100011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110100011000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110100011000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110100011000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110100011000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110100011000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100011001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110100011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110100011001010) && ({row_reg, col_reg}<19'b0111110100011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100011011011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110100011011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110100011011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100011011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110100011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100011100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111110100011100001) && ({row_reg, col_reg}<19'b0111110100011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100011100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110100011100100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110100011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100011100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110100011100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100011101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110100011101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110100011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100011101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111110100011101100) && ({row_reg, col_reg}<19'b0111110100011101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100011101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110100011110000) && ({row_reg, col_reg}<19'b0111110100011110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110100011110011) && ({row_reg, col_reg}<19'b0111110100011110101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110100011110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111110100011110110) && ({row_reg, col_reg}<19'b0111110100011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110100011111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110100011111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110100011111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110100011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100011111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110100011111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110100011111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110100011111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100100000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110100100000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100100000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110100100000011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110100100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100100000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100100000110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111110100100000111) && ({row_reg, col_reg}<19'b0111110100100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110100100001001) && ({row_reg, col_reg}<19'b0111110100100001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110100100001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100100001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110100100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100100001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110100100001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110100100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110100100010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110100100010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110100100010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111110100100010100) && ({row_reg, col_reg}<19'b0111110100100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110100100100011) && ({row_reg, col_reg}<19'b0111110100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100100100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100100100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110100100101000) && ({row_reg, col_reg}<19'b0111110100100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110100100101010) && ({row_reg, col_reg}<19'b0111110100100101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110100100101100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111110100100101101) && ({row_reg, col_reg}<19'b0111110100100110000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110100100110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110100100110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100100110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111110100100110011) && ({row_reg, col_reg}<19'b0111110100100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110100100111000) && ({row_reg, col_reg}<19'b0111110100101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100101000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110100101000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111110100101000010) && ({row_reg, col_reg}<19'b0111110100101000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110100101000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111110100101000101) && ({row_reg, col_reg}<19'b0111110100101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100101000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100101001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110100101001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110100101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100101001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100101001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110100101001110) && ({row_reg, col_reg}<19'b0111110100101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100101010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110100101010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110100101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100101010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110100101010101) && ({row_reg, col_reg}<19'b0111110100101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110100101101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110100101101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111110100101101100) && ({row_reg, col_reg}<19'b0111110100101101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100101101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110100101101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110100101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110100101110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110100101110010) && ({row_reg, col_reg}<19'b0111110100101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100101110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110100101110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111110100101110110) && ({row_reg, col_reg}<19'b0111110100101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100101111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111110100101111001) && ({row_reg, col_reg}<19'b0111110100101111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100101111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111110100101111100) && ({row_reg, col_reg}<19'b0111110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100101111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100101111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111110100110000000) && ({row_reg, col_reg}<19'b0111110100110000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111110100110000010) && ({row_reg, col_reg}<19'b0111110100110000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100110000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110100110000101) && ({row_reg, col_reg}<19'b0111110100110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110100110001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110100110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100110001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110100110001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111110100110001101) && ({row_reg, col_reg}<19'b0111110100110001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0111110100110001111) && ({row_reg, col_reg}<19'b0111110100110010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110100110010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100110010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110100110010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110100110010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100110010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110100110010111) && ({row_reg, col_reg}<19'b0111110100110011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110100110011100) && ({row_reg, col_reg}<19'b0111110100110100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110100110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110100110100001) && ({row_reg, col_reg}<19'b0111110100110101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111110100110101000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111110100110101001)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0111110100110101010)) color_data = 12'b110110111101;
		if(({row_reg, col_reg}==19'b0111110100110101011)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0111110100110101100)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}==19'b0111110100110101101)) color_data = 12'b110010011100;
		if(({row_reg, col_reg}==19'b0111110100110101110)) color_data = 12'b101110001010;
		if(({row_reg, col_reg}==19'b0111110100110101111)) color_data = 12'b011101000110;
		if(({row_reg, col_reg}==19'b0111110100110110000)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111110100110110001)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111110100110110010)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==19'b0111110100110110011)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==19'b0111110100110110100)) color_data = 12'b111011001110;
		if(({row_reg, col_reg}==19'b0111110100110110101)) color_data = 12'b111011001101;
		if(({row_reg, col_reg}==19'b0111110100110110110)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==19'b0111110100110110111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==19'b0111110100110111000)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==19'b0111110100110111001)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}>=19'b0111110100110111010) && ({row_reg, col_reg}<19'b0111110100110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111110100110111111) && ({row_reg, col_reg}<19'b0111110101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110101001010001) && ({row_reg, col_reg}<19'b0111110101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111110101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111110101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111110110000000000) && ({row_reg, col_reg}<19'b0111110110010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110110010101010) && ({row_reg, col_reg}<19'b0111110110010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110110010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111110110010101110) && ({row_reg, col_reg}<19'b0111110110010110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110110010110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110110010110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110110010110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110010110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110010110101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110110010110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111110110010110111) && ({row_reg, col_reg}<19'b0111110110010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110110010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110110010111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110110010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110010111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110110011000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110011000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110011000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110110011000100) && ({row_reg, col_reg}<19'b0111110110011001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110011001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110110011001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111110110011001010) && ({row_reg, col_reg}<19'b0111110110011001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110110011001110) && ({row_reg, col_reg}<19'b0111110110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110011011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110110011011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110110011011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110110011100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110011100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111110110011100010) && ({row_reg, col_reg}<19'b0111110110011100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110011100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110110011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110011100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111110110011100111) && ({row_reg, col_reg}<19'b0111110110011101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110110011101001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110110011101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110110011101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110011101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110011101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110011101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110110011101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110110011110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110011110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110011110011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110011110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110011110101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111110110011110110) && ({row_reg, col_reg}<19'b0111110110011111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110110011111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110011111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110110011111010) && ({row_reg, col_reg}<19'b0111110110011111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110011111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110011111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110110011111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110110011111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110100000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110100000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110110100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110100000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110110100000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110110100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110110100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110100001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110110100001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110100001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110100001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111110110100001100) && ({row_reg, col_reg}<19'b0111110110100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110100001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111110110100001111) && ({row_reg, col_reg}<19'b0111110110100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110100010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110110100010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110100010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110100010100) && ({row_reg, col_reg}<19'b0111110110100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110110100100011) && ({row_reg, col_reg}<19'b0111110110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110100100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110110100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110100100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110100101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110110100101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110100101010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110110100101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111110110100101100) && ({row_reg, col_reg}<19'b0111110110100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110110100110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110100110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110100110011) && ({row_reg, col_reg}<19'b0111110110100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110110100111000) && ({row_reg, col_reg}<19'b0111110110101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110101000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110110101000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111110110101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110101000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110101000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110110101000101) && ({row_reg, col_reg}<19'b0111110110101000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110101000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110110101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110110101001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110110101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110101001101) && ({row_reg, col_reg}<19'b0111110110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110110101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110101010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110110101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110101010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110110101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111110110101010101) && ({row_reg, col_reg}<19'b0111110110101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110101101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110110101101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110110101101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111110110101101110) && ({row_reg, col_reg}<19'b0111110110101110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110101110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110110101110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111110110101110010) && ({row_reg, col_reg}<19'b0111110110101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111110110101110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110101110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110110101110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110101111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110101111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111110110101111011) && ({row_reg, col_reg}<19'b0111110110101111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110110101111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110110101111111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110110110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110110000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110110000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110110000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110110110000100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111110110110000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110110000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110110000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110110110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110110001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110110110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110110001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110110001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110110110001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110110001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110110001111) && ({row_reg, col_reg}<19'b0111110110110010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110110110010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110110110010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111110110110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111110110110010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111110110110010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110110010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111110110110010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111110110110011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111110110110011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111110110110011010) && ({row_reg, col_reg}<19'b0111110110110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110110110100001) && ({row_reg, col_reg}<19'b0111110110110101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111110110110101001)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==19'b0111110110110101010)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==19'b0111110110110101011)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==19'b0111110110110101100)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==19'b0111110110110101101)) color_data = 12'b011101000110;
		if(({row_reg, col_reg}==19'b0111110110110101110)) color_data = 12'b011000110101;
		if(({row_reg, col_reg}>=19'b0111110110110101111) && ({row_reg, col_reg}<19'b0111110110110110001)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111110110110110001)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111110110110110010)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==19'b0111110110110110011)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==19'b0111110110110110100)) color_data = 12'b111010111101;
		if(({row_reg, col_reg}==19'b0111110110110110101)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==19'b0111110110110110110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==19'b0111110110110110111)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==19'b0111110110110111000)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=19'b0111110110110111001) && ({row_reg, col_reg}<19'b0111110110110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111110110110111111) && ({row_reg, col_reg}<19'b0111110111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111110111001010001) && ({row_reg, col_reg}<19'b0111110111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111110111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111110111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111111000000000000) && ({row_reg, col_reg}<19'b0111111000010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111000010101010) && ({row_reg, col_reg}<19'b0111111000010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111000010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111111000010101110) && ({row_reg, col_reg}<19'b0111111000010110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000010110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111000010110110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111111000010110111) && ({row_reg, col_reg}<19'b0111111000010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000010111001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111000010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111000010111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111000010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111000010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111000010111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111000010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000011000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111000011000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111000011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000011000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111000011000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000011000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111111000011000111) && ({row_reg, col_reg}<19'b0111111000011001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111000011001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111000011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111000011001011) && ({row_reg, col_reg}<19'b0111111000011001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111000011001110) && ({row_reg, col_reg}<19'b0111111000011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111000011011001) && ({row_reg, col_reg}<19'b0111111000011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111000011011100) && ({row_reg, col_reg}<19'b0111111000011011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111000011011110) && ({row_reg, col_reg}<19'b0111111000011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000011100001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111000011100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000011100100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111111000011100101) && ({row_reg, col_reg}<19'b0111111000011100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111000011100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000011101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111000011101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111000011101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111000011101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111000011101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000011101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111000011101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111000011110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000011110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111000011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000011110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111000011110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000011110101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000011110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111000011110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111000011111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111000011111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111000011111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111000011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000011111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111000011111101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111000011111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111000011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111000100000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111000100000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111111000100000011) && ({row_reg, col_reg}<19'b0111111000100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111000100001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111111000100001010) && ({row_reg, col_reg}<19'b0111111000100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000100001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000100001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111000100001111) && ({row_reg, col_reg}<19'b0111111000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000100010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000100010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000100010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111000100010100) && ({row_reg, col_reg}<19'b0111111000100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111000100100011) && ({row_reg, col_reg}<19'b0111111000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000100100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111000100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000100100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111111000100101000) && ({row_reg, col_reg}<19'b0111111000100101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0111111000100101110) && ({row_reg, col_reg}<19'b0111111000100110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111000100110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111000100110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000100110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111000100110011) && ({row_reg, col_reg}<19'b0111111000100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111000100111000) && ({row_reg, col_reg}<19'b0111111000101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000101000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111000101000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111000101000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111000101000011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111000101000100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111000101000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111111000101000110) && ({row_reg, col_reg}<19'b0111111000101001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111111000101001000) && ({row_reg, col_reg}<19'b0111111000101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000101001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111000101001101) && ({row_reg, col_reg}<19'b0111111000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000101001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111000101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111000101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000101010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000101010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111111000101010101) && ({row_reg, col_reg}<19'b0111111000101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111000101101001) && ({row_reg, col_reg}<19'b0111111000101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000101101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111000101101110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111111000101101111) && ({row_reg, col_reg}<19'b0111111000101110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000101110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111000101110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111111000101110011) && ({row_reg, col_reg}<19'b0111111000101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111000101110101) && ({row_reg, col_reg}<19'b0111111000101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111000101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111000101111000) && ({row_reg, col_reg}<19'b0111111000101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000101111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111111000101111011) && ({row_reg, col_reg}<19'b0111111000101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000101111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111000101111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111000110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111000110000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111000110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111000110000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111000110000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000110000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111000110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000110001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000110001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111000110001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111000110001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111000110001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111000110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111000110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111000110010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000110010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000110010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111000110010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111111000110010101) && ({row_reg, col_reg}<19'b0111111000110010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000110010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111000110011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111000110011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111000110011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111000110011011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111000110011100) && ({row_reg, col_reg}<19'b0111111000110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111000110011110) && ({row_reg, col_reg}<19'b0111111000110100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111000110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111000110100001) && ({row_reg, col_reg}<19'b0111111000110101001)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111111000110101001)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111111000110101010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111111000110101011)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111111000110101100)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111111000110101101)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111111000110101110)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111111000110101111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111111000110110000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111111000110110001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111111000110110010)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111111000110110011)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==19'b0111111000110110100)) color_data = 12'b011101000110;
		if(({row_reg, col_reg}==19'b0111111000110110101)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==19'b0111111000110110110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0111111000110110111)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0111111000110111000) && ({row_reg, col_reg}<19'b0111111000110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111111000110111111) && ({row_reg, col_reg}<19'b0111111001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111001001010001) && ({row_reg, col_reg}<19'b0111111001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111111001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111111001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111111010000000000) && ({row_reg, col_reg}<19'b0111111010010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111010010101010) && ({row_reg, col_reg}<19'b0111111010010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111010010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111111010010101110) && ({row_reg, col_reg}<19'b0111111010010110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010010110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010010110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111010010110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111010010110100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111010010110101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111010010110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111010010110111) && ({row_reg, col_reg}<19'b0111111010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111010010111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111010010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111010010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111010010111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111010010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010011000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111010011000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010011000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111010011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111010011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010011000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111010011001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010011001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111010011001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111111010011001011) && ({row_reg, col_reg}<19'b0111111010011001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010011001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111010011001110) && ({row_reg, col_reg}<19'b0111111010011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111010011011001) && ({row_reg, col_reg}<19'b0111111010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010011011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111010011011110) && ({row_reg, col_reg}<19'b0111111010011100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111010011100000) && ({row_reg, col_reg}<19'b0111111010011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010011100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111010011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010011100100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010011100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111010011100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111010011100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010011101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010011101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010011101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111010011101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111010011101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010011101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111111010011101111) && ({row_reg, col_reg}<19'b0111111010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010011110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111010011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010011110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010011110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111010011110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111111010011110110) && ({row_reg, col_reg}<19'b0111111010011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010011111000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111010011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111010011111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111010011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010011111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111010011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111010011111110) && ({row_reg, col_reg}<19'b0111111010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010100000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111010100000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111010100000011) && ({row_reg, col_reg}<19'b0111111010100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010100000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111010100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010100001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111111010100001010) && ({row_reg, col_reg}<19'b0111111010100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010100001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111010100001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111111010100001110) && ({row_reg, col_reg}<19'b0111111010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111010100010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111010100010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010100010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111111010100010100) && ({row_reg, col_reg}<19'b0111111010100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010100010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111010100010111) && ({row_reg, col_reg}<19'b0111111010100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111010100100011) && ({row_reg, col_reg}<19'b0111111010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010100100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111010100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010100100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111010100101000) && ({row_reg, col_reg}<19'b0111111010100101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111010100101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111010100101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111010100101100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111010100101101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111010100101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111010100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111010100110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111010100110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010100110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111111010100110011) && ({row_reg, col_reg}<19'b0111111010100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111010100111000) && ({row_reg, col_reg}<19'b0111111010101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111010101000001) && ({row_reg, col_reg}<19'b0111111010101000011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111111010101000011) && ({row_reg, col_reg}<19'b0111111010101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010101000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111010101000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111010101001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111010101001101) && ({row_reg, col_reg}<19'b0111111010101010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010101010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111010101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010101010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111010101010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111111010101010101) && ({row_reg, col_reg}<19'b0111111010101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111010101101000) && ({row_reg, col_reg}<19'b0111111010101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111010101101010) && ({row_reg, col_reg}<19'b0111111010101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010101101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111010101101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111111010101110000) && ({row_reg, col_reg}<19'b0111111010101110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010101110010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111010101110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111010101110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111010101110101) && ({row_reg, col_reg}<19'b0111111010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010101111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010101111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111010101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111010101111100) && ({row_reg, col_reg}<19'b0111111010101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010101111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111010101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010110000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111010110000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111010110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010110000011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111010110000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111111010110000101) && ({row_reg, col_reg}<19'b0111111010110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010110000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111010110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010110001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111010110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010110001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111010110001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010110001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111010110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111010110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111010110010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111010110010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0111111010110010010) && ({row_reg, col_reg}<19'b0111111010110010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010110010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111010110011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010110011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010110011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111010110011011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111010110011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111010110011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111010110011110) && ({row_reg, col_reg}<19'b0111111010110100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111010110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111010110100001) && ({row_reg, col_reg}<19'b0111111010110101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111111010110101000)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==19'b0111111010110101001)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0111111010110101010) && ({row_reg, col_reg}<19'b0111111010110101110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111111010110101110) && ({row_reg, col_reg}<19'b0111111010110110000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111111010110110000)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}>=19'b0111111010110110001) && ({row_reg, col_reg}<19'b0111111010110110011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111111010110110011)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111111010110110100)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111111010110110101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0111111010110110110) && ({row_reg, col_reg}<19'b0111111010110111000)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111111010110111000) && ({row_reg, col_reg}<19'b0111111010111000000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}>=19'b0111111010111000000) && ({row_reg, col_reg}<19'b0111111011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111011001010001) && ({row_reg, col_reg}<19'b0111111011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111111011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111111011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111111100000000000) && ({row_reg, col_reg}<19'b0111111100010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111100010101010) && ({row_reg, col_reg}<19'b0111111100010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111111100010101110) && ({row_reg, col_reg}<19'b0111111100010110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100010110000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111100010110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111100010110010) && ({row_reg, col_reg}<19'b0111111100010110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100010110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111111100010111010) && ({row_reg, col_reg}<19'b0111111100010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111100010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100010111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111100010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100011000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111100011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111100011000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111100011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100011000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0111111100011000101) && ({row_reg, col_reg}<19'b0111111100011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100011000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100011001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100011001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111100011001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111111100011001011) && ({row_reg, col_reg}<19'b0111111100011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100011011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100011011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111100011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100011100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111100011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100011100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111100011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100011100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111100011100111) && ({row_reg, col_reg}<19'b0111111100011101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111100011101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111100011101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100011101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111100011101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100011101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111100011101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111100011101111) && ({row_reg, col_reg}<19'b0111111100011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100011110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111100011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100011110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111100011110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111100011110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111111100011110110) && ({row_reg, col_reg}<19'b0111111100011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100011111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111100011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100011111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111100011111101) && ({row_reg, col_reg}<19'b0111111100011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100011111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111100100000000) && ({row_reg, col_reg}<19'b0111111100100000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111111100100000011) && ({row_reg, col_reg}<19'b0111111100100000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100100000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111100100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100100001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111111100100001010) && ({row_reg, col_reg}<19'b0111111100100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100100001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111100100001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111100100001111) && ({row_reg, col_reg}<19'b0111111100100010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111100100010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111100100010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100100010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111100100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111100100010111) && ({row_reg, col_reg}<19'b0111111100100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100100100010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111100100100011) && ({row_reg, col_reg}<19'b0111111100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111100100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100100100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111100100101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111100100101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111100100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111100100101011) && ({row_reg, col_reg}<19'b0111111100100110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111100100110000) && ({row_reg, col_reg}<19'b0111111100100110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100100110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111100100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111100100110100) && ({row_reg, col_reg}<19'b0111111100100110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111100100110110) && ({row_reg, col_reg}<19'b0111111100101000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111100101000001) && ({row_reg, col_reg}<19'b0111111100101000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111100101000011) && ({row_reg, col_reg}<19'b0111111100101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111100101000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111100101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100101001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111100101001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111100101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111100101001101) && ({row_reg, col_reg}<19'b0111111100101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100101010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111100101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100101010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111100101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111100101010101) && ({row_reg, col_reg}<19'b0111111100101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111100101101010) && ({row_reg, col_reg}<19'b0111111100101101100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111100101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111100101101101) && ({row_reg, col_reg}<19'b0111111100101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100101110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111100101110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111100101110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100101110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111100101110100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111111100101110101) && ({row_reg, col_reg}<19'b0111111100101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100101111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111100101111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111100101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111100101111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111100101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100101111110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111100101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100110000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111100110000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111100110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100110000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111100110000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111100110000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100110000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111100110000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111100110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100110001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111100110001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111100110001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111100110001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100110001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111100110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111100110001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111100110010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111100110010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111100110010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111100110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100110010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111100110010101) && ({row_reg, col_reg}<19'b0111111100110010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111111100110010111) && ({row_reg, col_reg}<19'b0111111100110011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111100110011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111100110011010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111100110011011) && ({row_reg, col_reg}<19'b0111111100110100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111100110100001) && ({row_reg, col_reg}<19'b0111111100110101000)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111111100110101000)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111111100110101001)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}>=19'b0111111100110101010) && ({row_reg, col_reg}<19'b0111111100110101100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111111100110101100) && ({row_reg, col_reg}<19'b0111111100110101110)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0111111100110101110) && ({row_reg, col_reg}<19'b0111111100110110000)) color_data = 12'b001100000010;
		if(({row_reg, col_reg}==19'b0111111100110110000)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==19'b0111111100110110001)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111111100110110010)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111111100110110011)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==19'b0111111100110110100)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==19'b0111111100110110101)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111111100110110110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111111100110110111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=19'b0111111100110111000) && ({row_reg, col_reg}<19'b0111111100110111010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111111100110111010) && ({row_reg, col_reg}<19'b0111111100110111111)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111111100110111111)) color_data = 12'b000000010001;
		if(({row_reg, col_reg}>=19'b0111111100111000000) && ({row_reg, col_reg}<19'b0111111101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111101001010001) && ({row_reg, col_reg}<19'b0111111101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111111101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111111101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b0111111110000000000) && ({row_reg, col_reg}<19'b0111111110010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111110010101010) && ({row_reg, col_reg}<19'b0111111110010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111111110010101110) && ({row_reg, col_reg}<19'b0111111110010110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0111111110010110000) && ({row_reg, col_reg}<19'b0111111110010110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110010110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111110010110011) && ({row_reg, col_reg}<19'b0111111110010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110010111001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111111110010111010) && ({row_reg, col_reg}<19'b0111111110010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110010111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111110010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110010111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111110010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110011000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111110011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110011000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111110011000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111110011001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110011001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110011001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b0111111110011001011) && ({row_reg, col_reg}<19'b0111111110011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111111110011011010) && ({row_reg, col_reg}<19'b0111111110011011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111110011011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111111110011011101) && ({row_reg, col_reg}<19'b0111111110011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011100000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111110011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110011100100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0111111110011100101) && ({row_reg, col_reg}<19'b0111111110011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110011101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111110011101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110011101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111110011101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111111110011101110) && ({row_reg, col_reg}<19'b0111111110011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111110011110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111110011110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110011110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110011110101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110011110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111110011110111) && ({row_reg, col_reg}<19'b0111111110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111110011111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110011111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0111111110011111101) && ({row_reg, col_reg}<19'b0111111110011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110011111111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110100000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110100000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111110100000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b0111111110100000011) && ({row_reg, col_reg}<19'b0111111110100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110100000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111110100001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111110100001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0111111110100001010) && ({row_reg, col_reg}<19'b0111111110100001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111110100001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111110100001101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111110100001111) && ({row_reg, col_reg}<19'b0111111110100010001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111110100010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111110100010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0111111110100010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111110100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110100010101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111110100010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111111110100010111) && ({row_reg, col_reg}<19'b0111111110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110100100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111110100100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111110100101001) && ({row_reg, col_reg}<19'b0111111110100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110100101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111110100101110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111110100101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111110100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110100110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111110100110010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111110100110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110100110101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111110100110110) && ({row_reg, col_reg}<19'b0111111110101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110101000010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111110101000011) && ({row_reg, col_reg}<19'b0111111110101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110101000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110101000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111110101000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110101001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111110101001101) && ({row_reg, col_reg}<19'b0111111110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110101010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111110101010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110101010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111110101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111110101010101) && ({row_reg, col_reg}<19'b0111111110101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110101101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111110101101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b0111111110101101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b0111111110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111110101101111) && ({row_reg, col_reg}<19'b0111111110101110001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111110101110010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111110101110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110101110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b0111111110101110101) && ({row_reg, col_reg}<19'b0111111110101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110101111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0111111110101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111110101111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b0111111110101111100) && ({row_reg, col_reg}<19'b0111111110101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110101111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111110101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110110000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111111110110000001) && ({row_reg, col_reg}<19'b0111111110110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110110000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111110110000100) && ({row_reg, col_reg}<19'b0111111110110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110110000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111110110001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b0111111110110001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b0111111110110001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0111111110110001011) && ({row_reg, col_reg}<19'b0111111110110001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110110001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111110110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110110001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b0111111110110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111110110010001) && ({row_reg, col_reg}<19'b0111111110110010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b0111111110110010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b0111111110110010101) && ({row_reg, col_reg}<19'b0111111110110010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110110010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b0111111110110011000) && ({row_reg, col_reg}<19'b0111111110110101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110110101000)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==19'b0111111110110101001)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==19'b0111111110110101010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0111111110110101011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0111111110110101100) && ({row_reg, col_reg}<19'b0111111110110101110)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111111110110101110)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111111110110101111)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111111110110110000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=19'b0111111110110110001) && ({row_reg, col_reg}<19'b0111111110110110011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0111111110110110011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==19'b0111111110110110100)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==19'b0111111110110110101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==19'b0111111110110110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110110110111)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111111110110111000) && ({row_reg, col_reg}<19'b0111111110110111010)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==19'b0111111110110111010)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}>=19'b0111111110110111011) && ({row_reg, col_reg}<19'b0111111110110111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b0111111110110111110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111111110110111111)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}>=19'b0111111110111000000) && ({row_reg, col_reg}<19'b0111111111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b0111111111001010001) && ({row_reg, col_reg}<19'b0111111111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b0111111111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b0111111111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000000000000000000) && ({row_reg, col_reg}<19'b1000000000010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000000010101010) && ({row_reg, col_reg}<19'b1000000000010101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000000010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000010101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000010101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000010101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000000010110001) && ({row_reg, col_reg}<19'b1000000000010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000000010111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000000010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000010111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000000010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000011000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000000011000001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000000011000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000000011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000011000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1000000000011000101) && ({row_reg, col_reg}<19'b1000000000011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000011000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000000011001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000011001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000000011001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000000000011001011) && ({row_reg, col_reg}<19'b1000000000011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000011011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000000011011010) && ({row_reg, col_reg}<19'b1000000000011011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000011011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000011011110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000000011011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000000011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000011100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b1000000000011100010) && ({row_reg, col_reg}<19'b1000000000011100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000011100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b1000000000011100101) && ({row_reg, col_reg}<19'b1000000000011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000011100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000000011101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1000000000011101001) && ({row_reg, col_reg}<19'b1000000000011101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000000011101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000000011101100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000000011101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000000011101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1000000000011101111) && ({row_reg, col_reg}<19'b1000000000011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000011110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000000011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000000011110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000000011110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000011110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000000011110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000000011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000000011111000) && ({row_reg, col_reg}<19'b1000000000011111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000000011111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000000011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000011111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000000011111101) && ({row_reg, col_reg}<19'b1000000000011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000011111111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000000100000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000000100000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000100000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000000100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000000100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000100000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000000100000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000000100000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000000100001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000000100001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1000000000100001010) && ({row_reg, col_reg}<19'b1000000000100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000100001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b1000000000100001101) && ({row_reg, col_reg}<19'b1000000000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000100010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000000100010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000100010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000000100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000100010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000000100010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000000000100010111) && ({row_reg, col_reg}<19'b1000000000100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000000100100001) && ({row_reg, col_reg}<19'b1000000000100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000000100100011) && ({row_reg, col_reg}<19'b1000000000100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000100100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000000100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000100101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000000100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000100101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000000100101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000000100101100) && ({row_reg, col_reg}<19'b1000000000100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000100101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000000100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000100110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000000100110010) && ({row_reg, col_reg}<19'b1000000000100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000100110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000000100111000) && ({row_reg, col_reg}<19'b1000000000101000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000101000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000000101000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000000101000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000000101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b1000000000101001000) && ({row_reg, col_reg}<19'b1000000000101001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000000101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000000101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000101001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1000000000101001101) && ({row_reg, col_reg}<19'b1000000000101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000000101010001) && ({row_reg, col_reg}<19'b1000000000101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000101010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b1000000000101010100) && ({row_reg, col_reg}<19'b1000000000101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000101010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000000101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000000101011000) && ({row_reg, col_reg}<19'b1000000000101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000101101001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000000101101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000000101101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000000101101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1000000000101101101) && ({row_reg, col_reg}<19'b1000000000101101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000101101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000000101110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000101110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000000101110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000101110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000000101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000000101110101) && ({row_reg, col_reg}<19'b1000000000101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000000101111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000000101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000000101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000000101111100) && ({row_reg, col_reg}<19'b1000000000101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000101111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000000101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000110000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000000110000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000000110000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000000110000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1000000000110000100) && ({row_reg, col_reg}<19'b1000000000110000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000110000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000000110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000110001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000110001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000000110001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000000110001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000000110001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000000110001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b1000000000110001110) && ({row_reg, col_reg}<19'b1000000000110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000000110010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000000110010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000000110010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000110010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000000000110011000) && ({row_reg, col_reg}<19'b1000000001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000001001010001) && ({row_reg, col_reg}<19'b1000000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000000001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000000001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000000010000000000) && ({row_reg, col_reg}<19'b1000000010010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010010101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000010010101001) && ({row_reg, col_reg}<19'b1000000010010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010010101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010010101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010010101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000010010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000010010110001) && ({row_reg, col_reg}<19'b1000000010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010010111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000010010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010010111100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000010010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010010111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000010010111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010011000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010011000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000010011000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010011000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000010011000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000010011000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000010011001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010011001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000010011001010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000010011001011) && ({row_reg, col_reg}<19'b1000000010011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010011011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000010011011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000010011011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000010011011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010011011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1000000010011011101) && ({row_reg, col_reg}<19'b1000000010011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010011011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000010011100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000010011100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010011100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010011100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010011100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b1000000010011100101) && ({row_reg, col_reg}<19'b1000000010011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010011100111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000010011101000) && ({row_reg, col_reg}<19'b1000000010011101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010011101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010011101011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000010011101100) && ({row_reg, col_reg}<19'b1000000010011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010011101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1000000010011101111) && ({row_reg, col_reg}<19'b1000000010011110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010011110001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010011110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000010011110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010011110100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010011110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000010011110110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000000010011110111) && ({row_reg, col_reg}<19'b1000000010011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000010011111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010011111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000010011111101) && ({row_reg, col_reg}<19'b1000000010100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000010100000001) && ({row_reg, col_reg}<19'b1000000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000010100000100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010100000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1000000010100000110) && ({row_reg, col_reg}<19'b1000000010100001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000010100001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000010100001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000010100001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010100001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010100001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000010100001101) && ({row_reg, col_reg}<19'b1000000010100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000010100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010100010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000010100010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010100010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000010100010100) && ({row_reg, col_reg}<19'b1000000010100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010100010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000010100010111) && ({row_reg, col_reg}<19'b1000000010100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000010100100001) && ({row_reg, col_reg}<19'b1000000010100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000010100100011) && ({row_reg, col_reg}<19'b1000000010100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010100100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010100100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010100101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000010100101001) && ({row_reg, col_reg}<19'b1000000010100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010100101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000010100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000010100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010100101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010100101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010100110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b1000000010100110010) && ({row_reg, col_reg}<19'b1000000010100110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010100110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000010100111000) && ({row_reg, col_reg}<19'b1000000010101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010101000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010101000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000010101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010101001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000010101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010101001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000010101001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000010101001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010101001110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000010101001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010101010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000010101010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010101010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000010101010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000010101010100) && ({row_reg, col_reg}<19'b1000000010101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010101010110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000010101010111) && ({row_reg, col_reg}<19'b1000000010101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010101101000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000010101101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000010101101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010101101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010101101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000010101101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010101101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000010101110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1000000010101110001) && ({row_reg, col_reg}<19'b1000000010101110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010101110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000010101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000010101110101) && ({row_reg, col_reg}<19'b1000000010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000010101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000010101111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010101111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000010101111100) && ({row_reg, col_reg}<19'b1000000010101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010101111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b1000000010101111111) && ({row_reg, col_reg}<19'b1000000010110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000010110000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000010110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010110000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1000000010110000101) && ({row_reg, col_reg}<19'b1000000010110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010110000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000010110001000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010110001001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000010110001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000010110001011) && ({row_reg, col_reg}<19'b1000000010110001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010110001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000010110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010110001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000010110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000010110010001) && ({row_reg, col_reg}<19'b1000000010110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000010110010100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000010110010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000010110010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010110010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000010110011000) && ({row_reg, col_reg}<19'b1000000011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000011001010001) && ({row_reg, col_reg}<19'b1000000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000000011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000000011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000000100000000000) && ({row_reg, col_reg}<19'b1000000100010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b1000000100010101110) && ({row_reg, col_reg}<19'b1000000100010110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000100010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000100010110001) && ({row_reg, col_reg}<19'b1000000100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000100010111010) && ({row_reg, col_reg}<19'b1000000100010111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100010111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000100010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000100010111111) && ({row_reg, col_reg}<19'b1000000100011000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100011000001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000100011000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000100011000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000100011000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100011000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100011000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000100011000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100011001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000100011001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000100011001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000100011001011) && ({row_reg, col_reg}<19'b1000000100011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000100011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100011011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b1000000100011011011) && ({row_reg, col_reg}<19'b1000000100011011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100011011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000100011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100011011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000100011100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000100011100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100011100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000100011100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000100011100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000000100011100101) && ({row_reg, col_reg}<19'b1000000100011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100011100111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000100011101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000100011101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000100011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000100011101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000100011101100) && ({row_reg, col_reg}<19'b1000000100011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100011101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000100011101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100011110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000100011110001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000100011110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100011110011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000100011110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000100011110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000100011110110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000100011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000100011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000100011111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000100011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100011111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000100011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000100011111110) && ({row_reg, col_reg}<19'b1000000100100000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100100000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1000000100100000010) && ({row_reg, col_reg}<19'b1000000100100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100100000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000100100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000100100001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000100100001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000100100001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000100100001101) && ({row_reg, col_reg}<19'b1000000100100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100100010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000100100010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100100010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000100100010100) && ({row_reg, col_reg}<19'b1000000100100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000100100010110) && ({row_reg, col_reg}<19'b1000000100100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000100100011000) && ({row_reg, col_reg}<19'b1000000100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100100100101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000100100100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000100100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000100100101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000100100101010) && ({row_reg, col_reg}<19'b1000000100100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100100101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000100100101110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100100101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100100110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000100100110001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000100100110010) && ({row_reg, col_reg}<19'b1000000100100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000100100110101) && ({row_reg, col_reg}<19'b1000000100101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100101000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000100101000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100101001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000100101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100101001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000100101001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1000000100101001100) && ({row_reg, col_reg}<19'b1000000100101001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100101001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000100101001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000100101010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100101010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100101010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000100101010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000100101010100) && ({row_reg, col_reg}<19'b1000000100101101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000100101101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000100101101011) && ({row_reg, col_reg}<19'b1000000100101101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100101101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100101101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000100101101111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000100101110000) && ({row_reg, col_reg}<19'b1000000100101110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100101110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100101110011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000100101110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000100101110101) && ({row_reg, col_reg}<19'b1000000100101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000100101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100101111000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000100101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100101111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000100101111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000000100101111100) && ({row_reg, col_reg}<19'b1000000100101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100101111110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000100101111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000100110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100110000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1000000100110000010) && ({row_reg, col_reg}<19'b1000000100110000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1000000100110000100) && ({row_reg, col_reg}<19'b1000000100110000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000100110000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000100110000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100110001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000100110001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000100110001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000100110001011) && ({row_reg, col_reg}<19'b1000000100110001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100110001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000100110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100110001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000100110010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000100110010001) && ({row_reg, col_reg}<19'b1000000100110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000100110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000100110010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100110010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100110010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1000000100110011000) && ({row_reg, col_reg}<19'b1000000101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000101001010001) && ({row_reg, col_reg}<19'b1000000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000000101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000000101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000000110000000000) && ({row_reg, col_reg}<19'b1000000110010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110010101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000110010101110) && ({row_reg, col_reg}<19'b1000000110010110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000110010110001) && ({row_reg, col_reg}<19'b1000000110010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110010111001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000110010111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000110010111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110010111100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000110010111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000110010111111) && ({row_reg, col_reg}<19'b1000000110011000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000110011000001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000000110011000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000110011000011) && ({row_reg, col_reg}<19'b1000000110011000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110011000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000110011000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000110011001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000110011001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000110011001010) && ({row_reg, col_reg}<19'b1000000110011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000110011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110011011010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000110011011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000110011011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110011011101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000110011011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000110011011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000110011100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110011100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000110011100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000110011100011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000000110011100100) && ({row_reg, col_reg}<19'b1000000110011100111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000110011101000) && ({row_reg, col_reg}<19'b1000000110011101010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000110011101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000110011101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000110011101100) && ({row_reg, col_reg}<19'b1000000110011101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110011101111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110011110000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000110011110001) && ({row_reg, col_reg}<19'b1000000110011110011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110011110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000110011110101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000110011110110) && ({row_reg, col_reg}<19'b1000000110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110011111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110011111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000110011111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110011111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000110011111101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000110011111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000110011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110100000000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000110100000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000110100000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000110100000100) && ({row_reg, col_reg}<19'b1000000110100000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000110100000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000110100000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000110100001000) && ({row_reg, col_reg}<19'b1000000110100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000110100001010) && ({row_reg, col_reg}<19'b1000000110100001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000110100001100) && ({row_reg, col_reg}<19'b1000000110100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110100001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110100010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000110100010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000110100010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b1000000110100010100) && ({row_reg, col_reg}<19'b1000000110100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000110100010110) && ({row_reg, col_reg}<19'b1000000110100011000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000110100011000) && ({row_reg, col_reg}<19'b1000000110100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000110100100100) && ({row_reg, col_reg}<19'b1000000110100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000000110100101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000110100101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000110100101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110100101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110100101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1000000110100101110) && ({row_reg, col_reg}<19'b1000000110100110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110100110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000000110100110001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000110100110010) && ({row_reg, col_reg}<19'b1000000110100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000000110100110101) && ({row_reg, col_reg}<19'b1000000110101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110101000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000110101000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000110101000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000110101001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000110101001001) && ({row_reg, col_reg}<19'b1000000110101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110101001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1000000110101001101) && ({row_reg, col_reg}<19'b1000000110101010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110101010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000110101010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000110101010010) && ({row_reg, col_reg}<19'b1000000110101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000110101010101) && ({row_reg, col_reg}<19'b1000000110101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110101010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000000110101011000) && ({row_reg, col_reg}<19'b1000000110101101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110101101010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000000110101101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000110101101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1000000110101101101) && ({row_reg, col_reg}<19'b1000000110101110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110101110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1000000110101110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000110101110010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000110101110011) && ({row_reg, col_reg}<19'b1000000110101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000110101110101) && ({row_reg, col_reg}<19'b1000000110101110111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000110101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110101111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000110101111001) && ({row_reg, col_reg}<19'b1000000110101111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110101111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000000110101111100) && ({row_reg, col_reg}<19'b1000000110101111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110101111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000110101111111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000000110110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000110110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110110000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000110110000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000000110110000100) && ({row_reg, col_reg}<19'b1000000110110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110110000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110110000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000110110001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b1000000110110001001) && ({row_reg, col_reg}<19'b1000000110110001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110110001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000110110001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000110110001101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000000110110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110110001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000000110110010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000000110110010001) && ({row_reg, col_reg}<19'b1000000110110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000000110110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000110110010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000110110010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=19'b1000000110110011000) && ({row_reg, col_reg}<19'b1000000111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000000111001010001) && ({row_reg, col_reg}<19'b1000000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000000111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000000111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000001000000000000) && ({row_reg, col_reg}<19'b1000001000010101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000010101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000010101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1000001000010101110) && ({row_reg, col_reg}<19'b1000001000010110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000001000010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000010110001) && ({row_reg, col_reg}<19'b1000001000010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000010111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001000010111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000010111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000010111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001000010111110) && ({row_reg, col_reg}<19'b1000001000011000000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001000011000000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000001000011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000011000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000011000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000001000011000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001000011000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001000011000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000001000011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000011001000) && ({row_reg, col_reg}<19'b1000001000011011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000011011010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000011011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000001000011011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1000001000011011101) && ({row_reg, col_reg}<19'b1000001000011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001000011011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001000011100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001000011100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000001000011100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001000011100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001000011100100) && ({row_reg, col_reg}<19'b1000001000011100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000011100110) && ({row_reg, col_reg}<19'b1000001000011101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000011101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000011101101) && ({row_reg, col_reg}<19'b1000001000011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000011111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000001000011111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001000011111100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001000011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000011111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001000011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000100000001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001000100000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001000100000011) && ({row_reg, col_reg}<19'b1000001000100000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001000100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000100000111) && ({row_reg, col_reg}<19'b1000001000100010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000100010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001000100010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000001000100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001000100010101) && ({row_reg, col_reg}<19'b1000001000100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000100010111) && ({row_reg, col_reg}<19'b1000001000100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000100100000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001000100100001) && ({row_reg, col_reg}<19'b1000001000100100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000100100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001000100100100) && ({row_reg, col_reg}<19'b1000001000100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001000100100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1000001000100101000) && ({row_reg, col_reg}<19'b1000001000100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001000100101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001000100101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000100101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001000100101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001000100101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000001000100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001000100110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001000100110001) && ({row_reg, col_reg}<19'b1000001000100110100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000100110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000100110101) && ({row_reg, col_reg}<19'b1000001000101000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000101000101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000101000110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001000101000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000001000101001000) && ({row_reg, col_reg}<19'b1000001000101001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000101001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000101001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000001000101001101) && ({row_reg, col_reg}<19'b1000001000101001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000001000101001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000101010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000001000101010001) && ({row_reg, col_reg}<19'b1000001000101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000101010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000101010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001000101010101) && ({row_reg, col_reg}<19'b1000001000101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000101010111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001000101011000) && ({row_reg, col_reg}<19'b1000001000101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000101101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001000101101001) && ({row_reg, col_reg}<19'b1000001000101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000101101011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001000101101100) && ({row_reg, col_reg}<19'b1000001000101101111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001000101101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b1000001000101110000) && ({row_reg, col_reg}<19'b1000001000101110010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001000101110010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000101110011) && ({row_reg, col_reg}<19'b1000001000101110101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001000101110101) && ({row_reg, col_reg}<19'b1000001000101110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000101111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001000101111001) && ({row_reg, col_reg}<19'b1000001000101111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001000101111011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001000101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000101111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000101111110) && ({row_reg, col_reg}<19'b1000001000110000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000110000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000110000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000110000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001000110000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000110000100) && ({row_reg, col_reg}<19'b1000001000110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001000110000110) && ({row_reg, col_reg}<19'b1000001000110001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001000110001000) && ({row_reg, col_reg}<19'b1000001000110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001000110001100) && ({row_reg, col_reg}<19'b1000001000110001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001000110001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000110010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001000110010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000110010010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000110010011) && ({row_reg, col_reg}<19'b1000001000110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001000110010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001000110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000110010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001000110011000) && ({row_reg, col_reg}<19'b1000001001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001001001010001) && ({row_reg, col_reg}<19'b1000001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000001001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000001001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000001010000000000) && ({row_reg, col_reg}<19'b1000001010010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010010101010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010010101011) && ({row_reg, col_reg}<19'b1000001010010101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010010101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001010010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001010010101111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000001010010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010010110001) && ({row_reg, col_reg}<19'b1000001010010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010010111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001010010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001010010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001010010111100) && ({row_reg, col_reg}<19'b1000001010010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010010111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001010010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001010011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010011000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001010011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001010011000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001010011000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001010011000110) && ({row_reg, col_reg}<19'b1000001010011011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010011011001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010011011010) && ({row_reg, col_reg}<19'b1000001010011011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010011011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001010011011101) && ({row_reg, col_reg}<19'b1000001010011011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001010011011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000001010011100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001010011100001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010011100010) && ({row_reg, col_reg}<19'b1000001010011100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010011100101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010011100110) && ({row_reg, col_reg}<19'b1000001010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001010011101101) && ({row_reg, col_reg}<19'b1000001010011110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010011110000) && ({row_reg, col_reg}<19'b1000001010011110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010011110111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010011111000) && ({row_reg, col_reg}<19'b1000001010011111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010011111010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001010011111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001010011111100) && ({row_reg, col_reg}<19'b1000001010011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010011111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010011111111) && ({row_reg, col_reg}<19'b1000001010100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010100001001) && ({row_reg, col_reg}<19'b1000001010100010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001010100010101) && ({row_reg, col_reg}<19'b1000001010100010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010100010111) && ({row_reg, col_reg}<19'b1000001010100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001010100100000) && ({row_reg, col_reg}<19'b1000001010100100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010100100100) && ({row_reg, col_reg}<19'b1000001010100100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010100100110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001010100100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000001010100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001010100101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000001010100101010) && ({row_reg, col_reg}<19'b1000001010100101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001010100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001010100101111) && ({row_reg, col_reg}<19'b1000001010101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001010101001110) && ({row_reg, col_reg}<19'b1000001010101010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010101010000) && ({row_reg, col_reg}<19'b1000001010101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010101010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001010101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010101010101) && ({row_reg, col_reg}<19'b1000001010101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010101010111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010101011000) && ({row_reg, col_reg}<19'b1000001010101101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010101101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001010101101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010101101010) && ({row_reg, col_reg}<19'b1000001010101110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001010101110010) && ({row_reg, col_reg}<19'b1000001010101110100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001010101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010101110101) && ({row_reg, col_reg}<19'b1000001010101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010101111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001010101111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001010101111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001010101111011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001010101111100) && ({row_reg, col_reg}<19'b1000001010101111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010101111110) && ({row_reg, col_reg}<19'b1000001010110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010110000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001010110000100) && ({row_reg, col_reg}<19'b1000001010110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010110000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001010110000111) && ({row_reg, col_reg}<19'b1000001010110001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001010110001101) && ({row_reg, col_reg}<19'b1000001010110001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001010110001111) && ({row_reg, col_reg}<19'b1000001010110010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001010110010010) && ({row_reg, col_reg}<19'b1000001010110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001010110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001010110010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001010110010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001010110010111) && ({row_reg, col_reg}<19'b1000001011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001011001010001) && ({row_reg, col_reg}<19'b1000001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000001011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000001011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000001100000000000) && ({row_reg, col_reg}<19'b1000001100010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100010101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001100010101011) && ({row_reg, col_reg}<19'b1000001100010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100010101110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001100010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100010110001) && ({row_reg, col_reg}<19'b1000001100010111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100010111000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001100010111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001100010111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001100010111100) && ({row_reg, col_reg}<19'b1000001100010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100010111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001100010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001100011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100011000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001100011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001100011000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001100011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001100011000110) && ({row_reg, col_reg}<19'b1000001100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100011011101) && ({row_reg, col_reg}<19'b1000001100011011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001100011011111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100011100000) && ({row_reg, col_reg}<19'b1000001100011101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100011101000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001100011101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100011101010) && ({row_reg, col_reg}<19'b1000001100011101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100011101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001100011101111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001100011110000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100011110001) && ({row_reg, col_reg}<19'b1000001100011110011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100011110011) && ({row_reg, col_reg}<19'b1000001100011111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100011111011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100011111100) && ({row_reg, col_reg}<19'b1000001100011111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100011111110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001100011111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100100000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100100000001) && ({row_reg, col_reg}<19'b1000001100100000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100100000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001100100000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001100100001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100100001001) && ({row_reg, col_reg}<19'b1000001100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100100010001) && ({row_reg, col_reg}<19'b1000001100100100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100100100001) && ({row_reg, col_reg}<19'b1000001100100100011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100100100011) && ({row_reg, col_reg}<19'b1000001100100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100100100101) && ({row_reg, col_reg}<19'b1000001100100100111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001100100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100100101000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001100100101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100100101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001100100101011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001100100101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001100100101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100100101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001100100101111) && ({row_reg, col_reg}<19'b1000001100101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100101001001) && ({row_reg, col_reg}<19'b1000001100101001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001100101001011) && ({row_reg, col_reg}<19'b1000001100101001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100101001101) && ({row_reg, col_reg}<19'b1000001100101001111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100101001111) && ({row_reg, col_reg}<19'b1000001100101010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100101010011) && ({row_reg, col_reg}<19'b1000001100101010101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100101010101) && ({row_reg, col_reg}<19'b1000001100101101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100101101101) && ({row_reg, col_reg}<19'b1000001100101110000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001100101110000) && ({row_reg, col_reg}<19'b1000001100101110010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100101110010) && ({row_reg, col_reg}<19'b1000001100101110100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100101110100) && ({row_reg, col_reg}<19'b1000001100101110111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100101110111) && ({row_reg, col_reg}<19'b1000001100101111001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001100101111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000001100101111010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001100101111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001100101111101) && ({row_reg, col_reg}<19'b1000001100110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100110000010) && ({row_reg, col_reg}<19'b1000001100110000100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001100110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100110000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001100110000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=19'b1000001100110000111) && ({row_reg, col_reg}<19'b1000001100110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100110001110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001100110001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001100110010000) && ({row_reg, col_reg}<19'b1000001100110010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001100110010010) && ({row_reg, col_reg}<19'b1000001100110010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001100110010100) && ({row_reg, col_reg}<19'b1000001100110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001100110010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001100110010111) && ({row_reg, col_reg}<19'b1000001101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001101001010001) && ({row_reg, col_reg}<19'b1000001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000001101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000001101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000001110000000000) && ({row_reg, col_reg}<19'b1000001110010101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110010101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001110010101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110010101100) && ({row_reg, col_reg}<19'b1000001110010101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110010101110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001110010101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110010110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110010110001) && ({row_reg, col_reg}<19'b1000001110010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110010111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110010111011) && ({row_reg, col_reg}<19'b1000001110010111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110010111110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110010111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110011000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==19'b1000001110011000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001110011000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1000001110011000101) && ({row_reg, col_reg}<19'b1000001110011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110011001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001110011001001) && ({row_reg, col_reg}<19'b1000001110011001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110011001100) && ({row_reg, col_reg}<19'b1000001110011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110011011000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001110011011001) && ({row_reg, col_reg}<19'b1000001110011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001110011011011) && ({row_reg, col_reg}<19'b1000001110011011101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001110011011101) && ({row_reg, col_reg}<19'b1000001110011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110011011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001110011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001110011100001) && ({row_reg, col_reg}<19'b1000001110011100100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110011100100) && ({row_reg, col_reg}<19'b1000001110011101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001110011101001) && ({row_reg, col_reg}<19'b1000001110011101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110011101100) && ({row_reg, col_reg}<19'b1000001110011111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110011111000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110011111001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110011111010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110011111011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001110011111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110011111101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110011111110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001110011111111) && ({row_reg, col_reg}<19'b1000001110100000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110100000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110100000100) && ({row_reg, col_reg}<19'b1000001110100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110100001010)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110100001011) && ({row_reg, col_reg}<19'b1000001110100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110100010000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110100010001) && ({row_reg, col_reg}<19'b1000001110100010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110100010011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110100010100) && ({row_reg, col_reg}<19'b1000001110100010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110100010111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001110100011000) && ({row_reg, col_reg}<19'b1000001110100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110100100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001110100100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001110100100111) && ({row_reg, col_reg}<19'b1000001110100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110100101001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110100101010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001110100101011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110100101100) && ({row_reg, col_reg}<19'b1000001110100101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110100101111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001110100110000) && ({row_reg, col_reg}<19'b1000001110101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110101000001) && ({row_reg, col_reg}<19'b1000001110101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101001001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110101001010) && ({row_reg, col_reg}<19'b1000001110101001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001110101001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001110101001111) && ({row_reg, col_reg}<19'b1000001110101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110101010101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001110101010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001110101010111) && ({row_reg, col_reg}<19'b1000001110101101100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101101100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110101101101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001110101101110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110101101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101110000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110101110001) && ({row_reg, col_reg}<19'b1000001110101110110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101110110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110101110111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001110101111000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101111001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001110101111010) && ({row_reg, col_reg}<19'b1000001110101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101111100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110101111101) && ({row_reg, col_reg}<19'b1000001110101111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110101111111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001110110000000) && ({row_reg, col_reg}<19'b1000001110110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110110000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001110110000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000001110110000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110110000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000001110110000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==19'b1000001110110000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110110001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001110110001001) && ({row_reg, col_reg}<19'b1000001110110001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110110001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000001110110001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000001110110001101) && ({row_reg, col_reg}<19'b1000001110110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110110001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b1000001110110010000) && ({row_reg, col_reg}<19'b1000001110110010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001110110010010) && ({row_reg, col_reg}<19'b1000001110110010100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000001110110010100) && ({row_reg, col_reg}<19'b1000001110110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000001110110010110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000001110110010111) && ({row_reg, col_reg}<19'b1000001111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000001111001010001) && ({row_reg, col_reg}<19'b1000001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000001111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000001111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000010000000000000) && ({row_reg, col_reg}<19'b1000010000011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010000011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000010000011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010000011000010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=19'b1000010000011000011) && ({row_reg, col_reg}<19'b1000010000011000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010000011000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==19'b1000010000011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010000011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000010000011001000) && ({row_reg, col_reg}<19'b1000010001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000010001001010001) && ({row_reg, col_reg}<19'b1000010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000010001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000010001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000010010000000000) && ({row_reg, col_reg}<19'b1000010010011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010010011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000010010011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010010011000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b1000010010011000011) && ({row_reg, col_reg}<19'b1000010010011000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010010011000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000010010011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010010011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000010010011001000) && ({row_reg, col_reg}<19'b1000010011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000010011001010001) && ({row_reg, col_reg}<19'b1000010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000010011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000010011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000010100000000000) && ({row_reg, col_reg}<19'b1000010100011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010100011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000010100011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010100011000010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=19'b1000010100011000011) && ({row_reg, col_reg}<19'b1000010100011000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1000010100011000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==19'b1000010100011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010100011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000010100011001000) && ({row_reg, col_reg}<19'b1000010101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000010101001010001) && ({row_reg, col_reg}<19'b1000010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000010101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000010101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000010110000000000) && ({row_reg, col_reg}<19'b1000010110011000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000010110011000010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000010110011000011) && ({row_reg, col_reg}<19'b1000010110011000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010110011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000010110011000110) && ({row_reg, col_reg}<19'b1000010111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000010111001010001) && ({row_reg, col_reg}<19'b1000010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000010111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000010111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000011000000000000) && ({row_reg, col_reg}<19'b1000011000011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000011000011000000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000011000011000001) && ({row_reg, col_reg}<19'b1000011000011000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000011000011000011) && ({row_reg, col_reg}<19'b1000011000011000101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000011000011000101) && ({row_reg, col_reg}<19'b1000011000011000111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000011000011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000011000011001000) && ({row_reg, col_reg}<19'b1000011001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000011001001010001) && ({row_reg, col_reg}<19'b1000011001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000011001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000011001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000011010000000000) && ({row_reg, col_reg}<19'b1000011010011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000011010011000000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==19'b1000011010011000001)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000011010011000010) && ({row_reg, col_reg}<19'b1000011010011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==19'b1000011010011000110)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==19'b1000011010011000111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=19'b1000011010011001000) && ({row_reg, col_reg}<19'b1000011011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000011011001010001) && ({row_reg, col_reg}<19'b1000011011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000011011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000011011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000011100000000000) && ({row_reg, col_reg}<19'b1000011100011000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000011100011000000) && ({row_reg, col_reg}<19'b1000011100011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000011100011000011) && ({row_reg, col_reg}<19'b1000011100011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000011100011000101) && ({row_reg, col_reg}<19'b1000011100011001000)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000011100011001000) && ({row_reg, col_reg}<19'b1000011101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000011101001010001) && ({row_reg, col_reg}<19'b1000011101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000011101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000011101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000011110000000000) && ({row_reg, col_reg}<19'b1000011110011000001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000011110011000001) && ({row_reg, col_reg}<19'b1000011110011000011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000011110011000011) && ({row_reg, col_reg}<19'b1000011110011000101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000011110011000101) && ({row_reg, col_reg}<19'b1000011110011000111)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}>=19'b1000011110011000111) && ({row_reg, col_reg}<19'b1000011111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000011111001010001) && ({row_reg, col_reg}<19'b1000011111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000011111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000011111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000100000000000000) && ({row_reg, col_reg}<19'b1000100001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000100001001010001) && ({row_reg, col_reg}<19'b1000100001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000100001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000100001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000100010000000000) && ({row_reg, col_reg}<19'b1000100011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000100011001010001) && ({row_reg, col_reg}<19'b1000100011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000100011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000100011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000100100000000000) && ({row_reg, col_reg}<19'b1000100101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000100101001010001) && ({row_reg, col_reg}<19'b1000100101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000100101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000100101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000100110000000000) && ({row_reg, col_reg}<19'b1000100111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000100111001010001) && ({row_reg, col_reg}<19'b1000100111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000100111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000100111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000101000000000000) && ({row_reg, col_reg}<19'b1000101001001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000101001001010001) && ({row_reg, col_reg}<19'b1000101001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000101001001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000101001001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000101010000000000) && ({row_reg, col_reg}<19'b1000101011001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000101011001010001) && ({row_reg, col_reg}<19'b1000101011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000101011001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000101011001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000101100000000000) && ({row_reg, col_reg}<19'b1000101101001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000101101001010001) && ({row_reg, col_reg}<19'b1000101101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000101101001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000101101001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000101110000000000) && ({row_reg, col_reg}<19'b1000101111001010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000101111001010001) && ({row_reg, col_reg}<19'b1000101111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000101111001010110)) color_data = 12'b001000010011;

		if(({row_reg, col_reg}==19'b1000101111001010111)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}>=19'b1000110000000000000) && ({row_reg, col_reg}<19'b1000110001001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000110001001010000) && ({row_reg, col_reg}<19'b1000110001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000110001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1000110001001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1000110010000000000) && ({row_reg, col_reg}<19'b1000110011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000110011001010000) && ({row_reg, col_reg}<19'b1000110011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000110011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1000110011001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1000110100000000000) && ({row_reg, col_reg}<19'b1000110101001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000110101001010000) && ({row_reg, col_reg}<19'b1000110101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000110101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1000110101001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1000110110000000000) && ({row_reg, col_reg}<19'b1000110111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000110111001010000) && ({row_reg, col_reg}<19'b1000110111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000110111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1000110111001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1000111000000000000) && ({row_reg, col_reg}<19'b1000111001001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000111001001010000) && ({row_reg, col_reg}<19'b1000111001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000111001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1000111001001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1000111010000000000) && ({row_reg, col_reg}<19'b1000111011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000111011001010000) && ({row_reg, col_reg}<19'b1000111011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000111011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1000111011001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1000111100000000000) && ({row_reg, col_reg}<19'b1000111101001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000111101001010000) && ({row_reg, col_reg}<19'b1000111101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000111101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1000111101001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1000111110000000000) && ({row_reg, col_reg}<19'b1000111111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1000111111001010000) && ({row_reg, col_reg}<19'b1000111111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1000111111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1000111111001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001000000000000000) && ({row_reg, col_reg}<19'b1001000001001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001000001001010000) && ({row_reg, col_reg}<19'b1001000001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001000001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001000001001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001000010000000000) && ({row_reg, col_reg}<19'b1001000011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001000011001010000) && ({row_reg, col_reg}<19'b1001000011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001000011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001000011001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001000100000000000) && ({row_reg, col_reg}<19'b1001000101001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001000101001010000) && ({row_reg, col_reg}<19'b1001000101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001000101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001000101001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001000110000000000) && ({row_reg, col_reg}<19'b1001000111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001000111001010000) && ({row_reg, col_reg}<19'b1001000111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001000111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001000111001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001001000000000000) && ({row_reg, col_reg}<19'b1001001001001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001001001001010000) && ({row_reg, col_reg}<19'b1001001001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001001001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001001001001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001001010000000000) && ({row_reg, col_reg}<19'b1001001011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001001011001010000) && ({row_reg, col_reg}<19'b1001001011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001001011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001001011001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001001100000000000) && ({row_reg, col_reg}<19'b1001001101001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001001101001010000) && ({row_reg, col_reg}<19'b1001001101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001001101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001001101001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001001110000000000) && ({row_reg, col_reg}<19'b1001001111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001001111001010000) && ({row_reg, col_reg}<19'b1001001111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001001111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001001111001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001010000000000000) && ({row_reg, col_reg}<19'b1001010001001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001010001001010000) && ({row_reg, col_reg}<19'b1001010001001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001010001001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001010001001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001010010000000000) && ({row_reg, col_reg}<19'b1001010011001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001010011001010000) && ({row_reg, col_reg}<19'b1001010011001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001010011001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001010011001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001010100000000000) && ({row_reg, col_reg}<19'b1001010101001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001010101001010000) && ({row_reg, col_reg}<19'b1001010101001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001010101001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}==19'b1001010101001010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=19'b1001010110000000000) && ({row_reg, col_reg}<19'b1001010111001010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=19'b1001010111001010000) && ({row_reg, col_reg}<19'b1001010111001010110)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==19'b1001010111001010110)) color_data = 12'b000100010010;

		if(({row_reg, col_reg}>=19'b1001010111001010111) && ({row_reg, col_reg}<=19'b1001010111001010111)) color_data = 12'b001000100011;
	end
endmodule